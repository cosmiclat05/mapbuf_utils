module stencil_2d(
  // inputs
  input [31:0] orig_loadData,
  input [31:0] filter_loadData,
  input [31:0] sol_loadData,
  input  orig_start_valid,
  input  filter_start_valid,
  input  sol_start_valid,
  input  start_valid,
  input  clk,
  input  rst,
  input  out0_ready,
  input  orig_end_ready,
  input  filter_end_ready,
  input  sol_end_ready,
  input  end_ready,
  input  fork0_outs_0_valid__anchors_in,
  input  fork0_outs_0_ready__anchors_in,
  input  fork0_outs_1_valid__anchors_in,
  input  fork0_outs_1_ready__anchors_in,
  input  fork0_outs_2_valid__anchors_in,
  input  fork0_outs_2_ready__anchors_in,
  input  mem_controller0_memEnd_valid__anchors_in,
  input  mem_controller0_memEnd_ready__anchors_in,
  input [31:0] mem_controller1_ldData_0__data_anchors_in,
  input  mem_controller1_ldData_0_valid__anchors_in,
  input  mem_controller1_ldData_0_ready__anchors_in,
  input  mem_controller1_memEnd_valid__anchors_in,
  input  mem_controller1_memEnd_ready__anchors_in,
  input [31:0] mem_controller2_ldData_0__data_anchors_in,
  input  mem_controller2_ldData_0_valid__anchors_in,
  input  mem_controller2_ldData_0_ready__anchors_in,
  input  mem_controller2_memEnd_valid__anchors_in,
  input  mem_controller2_memEnd_ready__anchors_in,
  input  constant1_outs__data_anchors_in,
  input  constant1_outs_valid__anchors_in,
  input  constant1_outs_ready__anchors_in,
  input [5:0] extsi12_outs__data_anchors_in,
  input  extsi12_outs_valid__anchors_in,
  input  extsi12_outs_ready__anchors_in,
  input [5:0] buffer18_outs__data_anchors_in,
  input  buffer18_outs_valid__anchors_in,
  input  buffer18_outs_ready__anchors_in,
  input [5:0] buffer19_outs__data_anchors_in,
  input  buffer19_outs_valid__anchors_in,
  input  buffer19_outs_ready__anchors_in,
  input [5:0] mux8_outs__data_anchors_in,
  input  mux8_outs_valid__anchors_in,
  input  mux8_outs_ready__anchors_in,
  input  buffer20_outs_valid__anchors_in,
  input  buffer20_outs_ready__anchors_in,
  input  buffer21_outs_valid__anchors_in,
  input  buffer21_outs_ready__anchors_in,
  input  control_merge0_outs_valid__anchors_in,
  input  control_merge0_outs_ready__anchors_in,
  input  control_merge0_index__data_anchors_in,
  input  control_merge0_index_valid__anchors_in,
  input  control_merge0_index_ready__anchors_in,
  input  fork1_outs_0_valid__anchors_in,
  input  fork1_outs_0_ready__anchors_in,
  input  fork1_outs_1_valid__anchors_in,
  input  fork1_outs_1_ready__anchors_in,
  input  constant3_outs__data_anchors_in,
  input  constant3_outs_valid__anchors_in,
  input  constant3_outs_ready__anchors_in,
  input  fork2_outs_0__data_anchors_in,
  input  fork2_outs_0_valid__anchors_in,
  input  fork2_outs_0_ready__anchors_in,
  input  fork2_outs_1__data_anchors_in,
  input  fork2_outs_1_valid__anchors_in,
  input  fork2_outs_1_ready__anchors_in,
  input [2:0] extsi13_outs__data_anchors_in,
  input  extsi13_outs_valid__anchors_in,
  input  extsi13_outs_ready__anchors_in,
  input [31:0] extsi14_outs__data_anchors_in,
  input  extsi14_outs_valid__anchors_in,
  input  extsi14_outs_ready__anchors_in,
  input [2:0] buffer10_outs__data_anchors_in,
  input  buffer10_outs_valid__anchors_in,
  input  buffer10_outs_ready__anchors_in,
  input [2:0] buffer11_outs__data_anchors_in,
  input  buffer11_outs_valid__anchors_in,
  input  buffer11_outs_ready__anchors_in,
  input [2:0] mux9_outs__data_anchors_in,
  input  mux9_outs_valid__anchors_in,
  input  mux9_outs_ready__anchors_in,
  input [31:0] buffer12_outs__data_anchors_in,
  input  buffer12_outs_valid__anchors_in,
  input  buffer12_outs_ready__anchors_in,
  input [31:0] buffer13_outs__data_anchors_in,
  input  buffer13_outs_valid__anchors_in,
  input  buffer13_outs_ready__anchors_in,
  input [31:0] mux2_outs__data_anchors_in,
  input  mux2_outs_valid__anchors_in,
  input  mux2_outs_ready__anchors_in,
  input [5:0] buffer14_outs__data_anchors_in,
  input  buffer14_outs_valid__anchors_in,
  input  buffer14_outs_ready__anchors_in,
  input [5:0] buffer15_outs__data_anchors_in,
  input  buffer15_outs_valid__anchors_in,
  input  buffer15_outs_ready__anchors_in,
  input [5:0] mux10_outs__data_anchors_in,
  input  mux10_outs_valid__anchors_in,
  input  mux10_outs_ready__anchors_in,
  input  buffer16_outs_valid__anchors_in,
  input  buffer16_outs_ready__anchors_in,
  input  buffer17_outs_valid__anchors_in,
  input  buffer17_outs_ready__anchors_in,
  input  control_merge1_outs_valid__anchors_in,
  input  control_merge1_outs_ready__anchors_in,
  input  control_merge1_index__data_anchors_in,
  input  control_merge1_index_valid__anchors_in,
  input  control_merge1_index_ready__anchors_in,
  input  fork3_outs_0__data_anchors_in,
  input  fork3_outs_0_valid__anchors_in,
  input  fork3_outs_0_ready__anchors_in,
  input  fork3_outs_1__data_anchors_in,
  input  fork3_outs_1_valid__anchors_in,
  input  fork3_outs_1_ready__anchors_in,
  input  fork3_outs_2__data_anchors_in,
  input  fork3_outs_2_valid__anchors_in,
  input  fork3_outs_2_ready__anchors_in,
  input  fork4_outs_0_valid__anchors_in,
  input  fork4_outs_0_ready__anchors_in,
  input  fork4_outs_1_valid__anchors_in,
  input  fork4_outs_1_ready__anchors_in,
  input  constant4_outs__data_anchors_in,
  input  constant4_outs_valid__anchors_in,
  input  constant4_outs_ready__anchors_in,
  input [2:0] extsi15_outs__data_anchors_in,
  input  extsi15_outs_valid__anchors_in,
  input  extsi15_outs_ready__anchors_in,
  input [2:0] buffer0_outs__data_anchors_in,
  input  buffer0_outs_valid__anchors_in,
  input  buffer0_outs_ready__anchors_in,
  input [2:0] buffer1_outs__data_anchors_in,
  input  buffer1_outs_valid__anchors_in,
  input  buffer1_outs_ready__anchors_in,
  input [2:0] mux11_outs__data_anchors_in,
  input  mux11_outs_valid__anchors_in,
  input  mux11_outs_ready__anchors_in,
  input [2:0] fork5_outs_0__data_anchors_in,
  input  fork5_outs_0_valid__anchors_in,
  input  fork5_outs_0_ready__anchors_in,
  input [2:0] fork5_outs_1__data_anchors_in,
  input  fork5_outs_1_valid__anchors_in,
  input  fork5_outs_1_ready__anchors_in,
  input [2:0] fork5_outs_2__data_anchors_in,
  input  fork5_outs_2_valid__anchors_in,
  input  fork5_outs_2_ready__anchors_in,
  input [6:0] extsi16_outs__data_anchors_in,
  input  extsi16_outs_valid__anchors_in,
  input  extsi16_outs_ready__anchors_in,
  input [5:0] extsi17_outs__data_anchors_in,
  input  extsi17_outs_valid__anchors_in,
  input  extsi17_outs_ready__anchors_in,
  input [3:0] extsi18_outs__data_anchors_in,
  input  extsi18_outs_valid__anchors_in,
  input  extsi18_outs_ready__anchors_in,
  input [31:0] buffer2_outs__data_anchors_in,
  input  buffer2_outs_valid__anchors_in,
  input  buffer2_outs_ready__anchors_in,
  input [31:0] buffer3_outs__data_anchors_in,
  input  buffer3_outs_valid__anchors_in,
  input  buffer3_outs_ready__anchors_in,
  input [31:0] mux5_outs__data_anchors_in,
  input  mux5_outs_valid__anchors_in,
  input  mux5_outs_ready__anchors_in,
  input [5:0] buffer4_outs__data_anchors_in,
  input  buffer4_outs_valid__anchors_in,
  input  buffer4_outs_ready__anchors_in,
  input [5:0] buffer5_outs__data_anchors_in,
  input  buffer5_outs_valid__anchors_in,
  input  buffer5_outs_ready__anchors_in,
  input [5:0] mux12_outs__data_anchors_in,
  input  mux12_outs_valid__anchors_in,
  input  mux12_outs_ready__anchors_in,
  input [5:0] fork6_outs_0__data_anchors_in,
  input  fork6_outs_0_valid__anchors_in,
  input  fork6_outs_0_ready__anchors_in,
  input [5:0] fork6_outs_1__data_anchors_in,
  input  fork6_outs_1_valid__anchors_in,
  input  fork6_outs_1_ready__anchors_in,
  input [6:0] extsi19_outs__data_anchors_in,
  input  extsi19_outs_valid__anchors_in,
  input  extsi19_outs_ready__anchors_in,
  input [2:0] buffer6_outs__data_anchors_in,
  input  buffer6_outs_valid__anchors_in,
  input  buffer6_outs_ready__anchors_in,
  input [2:0] buffer7_outs__data_anchors_in,
  input  buffer7_outs_valid__anchors_in,
  input  buffer7_outs_ready__anchors_in,
  input [2:0] mux13_outs__data_anchors_in,
  input  mux13_outs_valid__anchors_in,
  input  mux13_outs_ready__anchors_in,
  input [2:0] fork7_outs_0__data_anchors_in,
  input  fork7_outs_0_valid__anchors_in,
  input  fork7_outs_0_ready__anchors_in,
  input [2:0] fork7_outs_1__data_anchors_in,
  input  fork7_outs_1_valid__anchors_in,
  input  fork7_outs_1_ready__anchors_in,
  input [2:0] fork7_outs_2__data_anchors_in,
  input  fork7_outs_2_valid__anchors_in,
  input  fork7_outs_2_ready__anchors_in,
  input [2:0] fork7_outs_3__data_anchors_in,
  input  fork7_outs_3_valid__anchors_in,
  input  fork7_outs_3_ready__anchors_in,
  input [8:0] extsi20_outs__data_anchors_in,
  input  extsi20_outs_valid__anchors_in,
  input  extsi20_outs_ready__anchors_in,
  input [4:0] extsi21_outs__data_anchors_in,
  input  extsi21_outs_valid__anchors_in,
  input  extsi21_outs_ready__anchors_in,
  input [3:0] extsi22_outs__data_anchors_in,
  input  extsi22_outs_valid__anchors_in,
  input  extsi22_outs_ready__anchors_in,
  input  buffer8_outs_valid__anchors_in,
  input  buffer8_outs_ready__anchors_in,
  input  buffer9_outs_valid__anchors_in,
  input  buffer9_outs_ready__anchors_in,
  input  control_merge2_outs_valid__anchors_in,
  input  control_merge2_outs_ready__anchors_in,
  input  control_merge2_index__data_anchors_in,
  input  control_merge2_index_valid__anchors_in,
  input  control_merge2_index_ready__anchors_in,
  input  fork8_outs_0__data_anchors_in,
  input  fork8_outs_0_valid__anchors_in,
  input  fork8_outs_0_ready__anchors_in,
  input  fork8_outs_1__data_anchors_in,
  input  fork8_outs_1_valid__anchors_in,
  input  fork8_outs_1_ready__anchors_in,
  input  fork8_outs_2__data_anchors_in,
  input  fork8_outs_2_valid__anchors_in,
  input  fork8_outs_2_ready__anchors_in,
  input  fork8_outs_3__data_anchors_in,
  input  fork8_outs_3_valid__anchors_in,
  input  fork8_outs_3_ready__anchors_in,
  input  source0_outs_valid__anchors_in,
  input  source0_outs_ready__anchors_in,
  input [5:0] constant5_outs__data_anchors_in,
  input  constant5_outs_valid__anchors_in,
  input  constant5_outs_ready__anchors_in,
  input [8:0] extsi23_outs__data_anchors_in,
  input  extsi23_outs_valid__anchors_in,
  input  extsi23_outs_ready__anchors_in,
  input  source1_outs_valid__anchors_in,
  input  source1_outs_ready__anchors_in,
  input [2:0] constant16_outs__data_anchors_in,
  input  constant16_outs_valid__anchors_in,
  input  constant16_outs_ready__anchors_in,
  input [3:0] extsi24_outs__data_anchors_in,
  input  extsi24_outs_valid__anchors_in,
  input  extsi24_outs_ready__anchors_in,
  input  source2_outs_valid__anchors_in,
  input  source2_outs_ready__anchors_in,
  input [1:0] constant17_outs__data_anchors_in,
  input  constant17_outs_valid__anchors_in,
  input  constant17_outs_ready__anchors_in,
  input [1:0] fork9_outs_0__data_anchors_in,
  input  fork9_outs_0_valid__anchors_in,
  input  fork9_outs_0_ready__anchors_in,
  input [1:0] fork9_outs_1__data_anchors_in,
  input  fork9_outs_1_valid__anchors_in,
  input  fork9_outs_1_ready__anchors_in,
  input [3:0] extui0_outs__data_anchors_in,
  input  extui0_outs_valid__anchors_in,
  input  extui0_outs_ready__anchors_in,
  input [3:0] extsi25_outs__data_anchors_in,
  input  extsi25_outs_valid__anchors_in,
  input  extsi25_outs_ready__anchors_in,
  input [3:0] shli1_result__data_anchors_in,
  input  shli1_result_valid__anchors_in,
  input  shli1_result_ready__anchors_in,
  input [4:0] extsi26_outs__data_anchors_in,
  input  extsi26_outs_valid__anchors_in,
  input  extsi26_outs_ready__anchors_in,
  input [4:0] addi8_result__data_anchors_in,
  input  addi8_result_valid__anchors_in,
  input  addi8_result_ready__anchors_in,
  input [5:0] extsi27_outs__data_anchors_in,
  input  extsi27_outs_valid__anchors_in,
  input  extsi27_outs_ready__anchors_in,
  input [5:0] addi9_result__data_anchors_in,
  input  addi9_result_valid__anchors_in,
  input  addi9_result_ready__anchors_in,
  input [31:0] extsi28_outs__data_anchors_in,
  input  extsi28_outs_valid__anchors_in,
  input  extsi28_outs_ready__anchors_in,
  input [31:0] mc_load0_addrOut__data_anchors_in,
  input  mc_load0_addrOut_valid__anchors_in,
  input  mc_load0_addrOut_ready__anchors_in,
  input [31:0] mc_load0_dataOut__data_anchors_in,
  input  mc_load0_dataOut_valid__anchors_in,
  input  mc_load0_dataOut_ready__anchors_in,
  input [6:0] addi10_result__data_anchors_in,
  input  addi10_result_valid__anchors_in,
  input  addi10_result_ready__anchors_in,
  input [9:0] extsi29_outs__data_anchors_in,
  input  extsi29_outs_valid__anchors_in,
  input  extsi29_outs_ready__anchors_in,
  input [8:0] muli1_result__data_anchors_in,
  input  muli1_result_valid__anchors_in,
  input  muli1_result_ready__anchors_in,
  input [9:0] extsi30_outs__data_anchors_in,
  input  extsi30_outs_valid__anchors_in,
  input  extsi30_outs_ready__anchors_in,
  input [9:0] addi11_result__data_anchors_in,
  input  addi11_result_valid__anchors_in,
  input  addi11_result_ready__anchors_in,
  input [31:0] extsi31_outs__data_anchors_in,
  input  extsi31_outs_valid__anchors_in,
  input  extsi31_outs_ready__anchors_in,
  input [31:0] mc_load1_addrOut__data_anchors_in,
  input  mc_load1_addrOut_valid__anchors_in,
  input  mc_load1_addrOut_ready__anchors_in,
  input [31:0] mc_load1_dataOut__data_anchors_in,
  input  mc_load1_dataOut_valid__anchors_in,
  input  mc_load1_dataOut_ready__anchors_in,
  input [31:0] muli0_result__data_anchors_in,
  input  muli0_result_valid__anchors_in,
  input  muli0_result_ready__anchors_in,
  input [31:0] addi0_result__data_anchors_in,
  input  addi0_result_valid__anchors_in,
  input  addi0_result_ready__anchors_in,
  input [3:0] addi12_result__data_anchors_in,
  input  addi12_result_valid__anchors_in,
  input  addi12_result_ready__anchors_in,
  input [3:0] fork10_outs_0__data_anchors_in,
  input  fork10_outs_0_valid__anchors_in,
  input  fork10_outs_0_ready__anchors_in,
  input [3:0] fork10_outs_1__data_anchors_in,
  input  fork10_outs_1_valid__anchors_in,
  input  fork10_outs_1_ready__anchors_in,
  input [2:0] trunci0_outs__data_anchors_in,
  input  trunci0_outs_valid__anchors_in,
  input  trunci0_outs_ready__anchors_in,
  input  cmpi3_result__data_anchors_in,
  input  cmpi3_result_valid__anchors_in,
  input  cmpi3_result_ready__anchors_in,
  input  fork11_outs_0__data_anchors_in,
  input  fork11_outs_0_valid__anchors_in,
  input  fork11_outs_0_ready__anchors_in,
  input  fork11_outs_1__data_anchors_in,
  input  fork11_outs_1_valid__anchors_in,
  input  fork11_outs_1_ready__anchors_in,
  input  fork11_outs_2__data_anchors_in,
  input  fork11_outs_2_valid__anchors_in,
  input  fork11_outs_2_ready__anchors_in,
  input  fork11_outs_3__data_anchors_in,
  input  fork11_outs_3_valid__anchors_in,
  input  fork11_outs_3_ready__anchors_in,
  input  fork11_outs_4__data_anchors_in,
  input  fork11_outs_4_valid__anchors_in,
  input  fork11_outs_4_ready__anchors_in,
  input [2:0] cond_br0_trueOut__data_anchors_in,
  input  cond_br0_trueOut_valid__anchors_in,
  input  cond_br0_trueOut_ready__anchors_in,
  input [2:0] cond_br0_falseOut__data_anchors_in,
  input  cond_br0_falseOut_valid__anchors_in,
  input  cond_br0_falseOut_ready__anchors_in,
  input [31:0] cond_br4_trueOut__data_anchors_in,
  input  cond_br4_trueOut_valid__anchors_in,
  input  cond_br4_trueOut_ready__anchors_in,
  input [31:0] cond_br4_falseOut__data_anchors_in,
  input  cond_br4_falseOut_valid__anchors_in,
  input  cond_br4_falseOut_ready__anchors_in,
  input [5:0] cond_br1_trueOut__data_anchors_in,
  input  cond_br1_trueOut_valid__anchors_in,
  input  cond_br1_trueOut_ready__anchors_in,
  input [5:0] cond_br1_falseOut__data_anchors_in,
  input  cond_br1_falseOut_valid__anchors_in,
  input  cond_br1_falseOut_ready__anchors_in,
  input [2:0] cond_br2_trueOut__data_anchors_in,
  input  cond_br2_trueOut_valid__anchors_in,
  input  cond_br2_trueOut_ready__anchors_in,
  input [2:0] cond_br2_falseOut__data_anchors_in,
  input  cond_br2_falseOut_valid__anchors_in,
  input  cond_br2_falseOut_ready__anchors_in,
  input  cond_br7_trueOut_valid__anchors_in,
  input  cond_br7_trueOut_ready__anchors_in,
  input  cond_br7_falseOut_valid__anchors_in,
  input  cond_br7_falseOut_ready__anchors_in,
  input [3:0] extsi32_outs__data_anchors_in,
  input  extsi32_outs_valid__anchors_in,
  input  extsi32_outs_ready__anchors_in,
  input  source3_outs_valid__anchors_in,
  input  source3_outs_ready__anchors_in,
  input [2:0] constant18_outs__data_anchors_in,
  input  constant18_outs_valid__anchors_in,
  input  constant18_outs_ready__anchors_in,
  input [3:0] extsi33_outs__data_anchors_in,
  input  extsi33_outs_valid__anchors_in,
  input  extsi33_outs_ready__anchors_in,
  input  source4_outs_valid__anchors_in,
  input  source4_outs_ready__anchors_in,
  input [1:0] constant19_outs__data_anchors_in,
  input  constant19_outs_valid__anchors_in,
  input  constant19_outs_ready__anchors_in,
  input [3:0] extsi34_outs__data_anchors_in,
  input  extsi34_outs_valid__anchors_in,
  input  extsi34_outs_ready__anchors_in,
  input [3:0] addi13_result__data_anchors_in,
  input  addi13_result_valid__anchors_in,
  input  addi13_result_ready__anchors_in,
  input [3:0] fork12_outs_0__data_anchors_in,
  input  fork12_outs_0_valid__anchors_in,
  input  fork12_outs_0_ready__anchors_in,
  input [3:0] fork12_outs_1__data_anchors_in,
  input  fork12_outs_1_valid__anchors_in,
  input  fork12_outs_1_ready__anchors_in,
  input [2:0] trunci1_outs__data_anchors_in,
  input  trunci1_outs_valid__anchors_in,
  input  trunci1_outs_ready__anchors_in,
  input  cmpi4_result__data_anchors_in,
  input  cmpi4_result_valid__anchors_in,
  input  cmpi4_result_ready__anchors_in,
  input  fork13_outs_0__data_anchors_in,
  input  fork13_outs_0_valid__anchors_in,
  input  fork13_outs_0_ready__anchors_in,
  input  fork13_outs_1__data_anchors_in,
  input  fork13_outs_1_valid__anchors_in,
  input  fork13_outs_1_ready__anchors_in,
  input  fork13_outs_2__data_anchors_in,
  input  fork13_outs_2_valid__anchors_in,
  input  fork13_outs_2_ready__anchors_in,
  input  fork13_outs_3__data_anchors_in,
  input  fork13_outs_3_valid__anchors_in,
  input  fork13_outs_3_ready__anchors_in,
  input [2:0] cond_br15_trueOut__data_anchors_in,
  input  cond_br15_trueOut_valid__anchors_in,
  input  cond_br15_trueOut_ready__anchors_in,
  input [2:0] cond_br15_falseOut__data_anchors_in,
  input  cond_br15_falseOut_valid__anchors_in,
  input  cond_br15_falseOut_ready__anchors_in,
  input [31:0] cond_br9_trueOut__data_anchors_in,
  input  cond_br9_trueOut_valid__anchors_in,
  input  cond_br9_trueOut_ready__anchors_in,
  input [31:0] cond_br9_falseOut__data_anchors_in,
  input  cond_br9_falseOut_valid__anchors_in,
  input  cond_br9_falseOut_ready__anchors_in,
  input [5:0] cond_br16_trueOut__data_anchors_in,
  input  cond_br16_trueOut_valid__anchors_in,
  input  cond_br16_trueOut_ready__anchors_in,
  input [5:0] cond_br16_falseOut__data_anchors_in,
  input  cond_br16_falseOut_valid__anchors_in,
  input  cond_br16_falseOut_ready__anchors_in,
  input  cond_br11_trueOut_valid__anchors_in,
  input  cond_br11_trueOut_ready__anchors_in,
  input  cond_br11_falseOut_valid__anchors_in,
  input  cond_br11_falseOut_ready__anchors_in,
  input [1:0] constant20_outs__data_anchors_in,
  input  constant20_outs_valid__anchors_in,
  input  constant20_outs_ready__anchors_in,
  input [31:0] extsi9_outs__data_anchors_in,
  input  extsi9_outs_valid__anchors_in,
  input  extsi9_outs_ready__anchors_in,
  input [5:0] fork14_outs_0__data_anchors_in,
  input  fork14_outs_0_valid__anchors_in,
  input  fork14_outs_0_ready__anchors_in,
  input [5:0] fork14_outs_1__data_anchors_in,
  input  fork14_outs_1_valid__anchors_in,
  input  fork14_outs_1_ready__anchors_in,
  input [6:0] extsi35_outs__data_anchors_in,
  input  extsi35_outs_valid__anchors_in,
  input  extsi35_outs_ready__anchors_in,
  input [31:0] extsi36_outs__data_anchors_in,
  input  extsi36_outs_valid__anchors_in,
  input  extsi36_outs_ready__anchors_in,
  input [31:0] fork15_outs_0__data_anchors_in,
  input  fork15_outs_0_valid__anchors_in,
  input  fork15_outs_0_ready__anchors_in,
  input [31:0] fork15_outs_1__data_anchors_in,
  input  fork15_outs_1_valid__anchors_in,
  input  fork15_outs_1_ready__anchors_in,
  input  fork16_outs_0_valid__anchors_in,
  input  fork16_outs_0_ready__anchors_in,
  input  fork16_outs_1_valid__anchors_in,
  input  fork16_outs_1_ready__anchors_in,
  input  source5_outs_valid__anchors_in,
  input  source5_outs_ready__anchors_in,
  input [5:0] constant21_outs__data_anchors_in,
  input  constant21_outs_valid__anchors_in,
  input  constant21_outs_ready__anchors_in,
  input [6:0] extsi37_outs__data_anchors_in,
  input  extsi37_outs_valid__anchors_in,
  input  extsi37_outs_ready__anchors_in,
  input  source6_outs_valid__anchors_in,
  input  source6_outs_ready__anchors_in,
  input [1:0] constant22_outs__data_anchors_in,
  input  constant22_outs_valid__anchors_in,
  input  constant22_outs_ready__anchors_in,
  input [6:0] extsi38_outs__data_anchors_in,
  input  extsi38_outs_valid__anchors_in,
  input  extsi38_outs_ready__anchors_in,
  input [31:0] mc_store0_addrOut__data_anchors_in,
  input  mc_store0_addrOut_valid__anchors_in,
  input  mc_store0_addrOut_ready__anchors_in,
  input [31:0] mc_store0_dataToMem__data_anchors_in,
  input  mc_store0_dataToMem_valid__anchors_in,
  input  mc_store0_dataToMem_ready__anchors_in,
  input [6:0] addi14_result__data_anchors_in,
  input  addi14_result_valid__anchors_in,
  input  addi14_result_ready__anchors_in,
  input [6:0] fork17_outs_0__data_anchors_in,
  input  fork17_outs_0_valid__anchors_in,
  input  fork17_outs_0_ready__anchors_in,
  input [6:0] fork17_outs_1__data_anchors_in,
  input  fork17_outs_1_valid__anchors_in,
  input  fork17_outs_1_ready__anchors_in,
  input [5:0] trunci2_outs__data_anchors_in,
  input  trunci2_outs_valid__anchors_in,
  input  trunci2_outs_ready__anchors_in,
  input  cmpi5_result__data_anchors_in,
  input  cmpi5_result_valid__anchors_in,
  input  cmpi5_result_ready__anchors_in,
  input  fork18_outs_0__data_anchors_in,
  input  fork18_outs_0_valid__anchors_in,
  input  fork18_outs_0_ready__anchors_in,
  input  fork18_outs_1__data_anchors_in,
  input  fork18_outs_1_valid__anchors_in,
  input  fork18_outs_1_ready__anchors_in,
  input  fork18_outs_2__data_anchors_in,
  input  fork18_outs_2_valid__anchors_in,
  input  fork18_outs_2_ready__anchors_in,
  input [5:0] cond_br17_trueOut__data_anchors_in,
  input  cond_br17_trueOut_valid__anchors_in,
  input  cond_br17_trueOut_ready__anchors_in,
  input [5:0] cond_br17_falseOut__data_anchors_in,
  input  cond_br17_falseOut_valid__anchors_in,
  input  cond_br17_falseOut_ready__anchors_in,
  input  cond_br13_trueOut_valid__anchors_in,
  input  cond_br13_trueOut_ready__anchors_in,
  input  cond_br13_falseOut_valid__anchors_in,
  input  cond_br13_falseOut_ready__anchors_in,
  input [31:0] cond_br14_trueOut__data_anchors_in,
  input  cond_br14_trueOut_valid__anchors_in,
  input  cond_br14_trueOut_ready__anchors_in,
  input [31:0] cond_br14_falseOut__data_anchors_in,
  input  cond_br14_falseOut_valid__anchors_in,
  input  cond_br14_falseOut_ready__anchors_in,
  input  fork19_outs_0_valid__anchors_in,
  input  fork19_outs_0_ready__anchors_in,
  input  fork19_outs_1_valid__anchors_in,
  input  fork19_outs_1_ready__anchors_in,
  input  fork19_outs_2_valid__anchors_in,
  input  fork19_outs_2_ready__anchors_in,
  // outputs
  output  orig_start_ready,
  output  filter_start_ready,
  output  sol_start_ready,
  output  start_ready,
  output [31:0] out0,
  output  out0_valid,
  output  orig_end_valid,
  output  filter_end_valid,
  output  sol_end_valid,
  output  end_valid,
  output  orig_loadEn,
  output [31:0] orig_loadAddr,
  output  orig_storeEn,
  output [31:0] orig_storeAddr,
  output [31:0] orig_storeData,
  output  filter_loadEn,
  output [31:0] filter_loadAddr,
  output  filter_storeEn,
  output [31:0] filter_storeAddr,
  output [31:0] filter_storeData,
  output  sol_loadEn,
  output [31:0] sol_loadAddr,
  output  sol_storeEn,
  output [31:0] sol_storeAddr,
  output [31:0] sol_storeData,
  output  fork0_outs_0_valid__anchors_out,
  output  fork0_outs_0_ready__anchors_out,
  output  fork0_outs_1_valid__anchors_out,
  output  fork0_outs_1_ready__anchors_out,
  output  fork0_outs_2_valid__anchors_out,
  output  fork0_outs_2_ready__anchors_out,
  output  mem_controller0_memEnd_valid__anchors_out,
  output  mem_controller0_memEnd_ready__anchors_out,
  output [31:0] mem_controller1_ldData_0__data_anchors_out,
  output  mem_controller1_ldData_0_valid__anchors_out,
  output  mem_controller1_ldData_0_ready__anchors_out,
  output  mem_controller1_memEnd_valid__anchors_out,
  output  mem_controller1_memEnd_ready__anchors_out,
  output [31:0] mem_controller2_ldData_0__data_anchors_out,
  output  mem_controller2_ldData_0_valid__anchors_out,
  output  mem_controller2_ldData_0_ready__anchors_out,
  output  mem_controller2_memEnd_valid__anchors_out,
  output  mem_controller2_memEnd_ready__anchors_out,
  output  constant1_outs__data_anchors_out,
  output  constant1_outs_valid__anchors_out,
  output  constant1_outs_ready__anchors_out,
  output [5:0] extsi12_outs__data_anchors_out,
  output  extsi12_outs_valid__anchors_out,
  output  extsi12_outs_ready__anchors_out,
  output [5:0] buffer18_outs__data_anchors_out,
  output  buffer18_outs_valid__anchors_out,
  output  buffer18_outs_ready__anchors_out,
  output [5:0] buffer19_outs__data_anchors_out,
  output  buffer19_outs_valid__anchors_out,
  output  buffer19_outs_ready__anchors_out,
  output [5:0] mux8_outs__data_anchors_out,
  output  mux8_outs_valid__anchors_out,
  output  mux8_outs_ready__anchors_out,
  output  buffer20_outs_valid__anchors_out,
  output  buffer20_outs_ready__anchors_out,
  output  buffer21_outs_valid__anchors_out,
  output  buffer21_outs_ready__anchors_out,
  output  control_merge0_outs_valid__anchors_out,
  output  control_merge0_outs_ready__anchors_out,
  output  control_merge0_index__data_anchors_out,
  output  control_merge0_index_valid__anchors_out,
  output  control_merge0_index_ready__anchors_out,
  output  fork1_outs_0_valid__anchors_out,
  output  fork1_outs_0_ready__anchors_out,
  output  fork1_outs_1_valid__anchors_out,
  output  fork1_outs_1_ready__anchors_out,
  output  constant3_outs__data_anchors_out,
  output  constant3_outs_valid__anchors_out,
  output  constant3_outs_ready__anchors_out,
  output  fork2_outs_0__data_anchors_out,
  output  fork2_outs_0_valid__anchors_out,
  output  fork2_outs_0_ready__anchors_out,
  output  fork2_outs_1__data_anchors_out,
  output  fork2_outs_1_valid__anchors_out,
  output  fork2_outs_1_ready__anchors_out,
  output [2:0] extsi13_outs__data_anchors_out,
  output  extsi13_outs_valid__anchors_out,
  output  extsi13_outs_ready__anchors_out,
  output [31:0] extsi14_outs__data_anchors_out,
  output  extsi14_outs_valid__anchors_out,
  output  extsi14_outs_ready__anchors_out,
  output [2:0] buffer10_outs__data_anchors_out,
  output  buffer10_outs_valid__anchors_out,
  output  buffer10_outs_ready__anchors_out,
  output [2:0] buffer11_outs__data_anchors_out,
  output  buffer11_outs_valid__anchors_out,
  output  buffer11_outs_ready__anchors_out,
  output [2:0] mux9_outs__data_anchors_out,
  output  mux9_outs_valid__anchors_out,
  output  mux9_outs_ready__anchors_out,
  output [31:0] buffer12_outs__data_anchors_out,
  output  buffer12_outs_valid__anchors_out,
  output  buffer12_outs_ready__anchors_out,
  output [31:0] buffer13_outs__data_anchors_out,
  output  buffer13_outs_valid__anchors_out,
  output  buffer13_outs_ready__anchors_out,
  output [31:0] mux2_outs__data_anchors_out,
  output  mux2_outs_valid__anchors_out,
  output  mux2_outs_ready__anchors_out,
  output [5:0] buffer14_outs__data_anchors_out,
  output  buffer14_outs_valid__anchors_out,
  output  buffer14_outs_ready__anchors_out,
  output [5:0] buffer15_outs__data_anchors_out,
  output  buffer15_outs_valid__anchors_out,
  output  buffer15_outs_ready__anchors_out,
  output [5:0] mux10_outs__data_anchors_out,
  output  mux10_outs_valid__anchors_out,
  output  mux10_outs_ready__anchors_out,
  output  buffer16_outs_valid__anchors_out,
  output  buffer16_outs_ready__anchors_out,
  output  buffer17_outs_valid__anchors_out,
  output  buffer17_outs_ready__anchors_out,
  output  control_merge1_outs_valid__anchors_out,
  output  control_merge1_outs_ready__anchors_out,
  output  control_merge1_index__data_anchors_out,
  output  control_merge1_index_valid__anchors_out,
  output  control_merge1_index_ready__anchors_out,
  output  fork3_outs_0__data_anchors_out,
  output  fork3_outs_0_valid__anchors_out,
  output  fork3_outs_0_ready__anchors_out,
  output  fork3_outs_1__data_anchors_out,
  output  fork3_outs_1_valid__anchors_out,
  output  fork3_outs_1_ready__anchors_out,
  output  fork3_outs_2__data_anchors_out,
  output  fork3_outs_2_valid__anchors_out,
  output  fork3_outs_2_ready__anchors_out,
  output  fork4_outs_0_valid__anchors_out,
  output  fork4_outs_0_ready__anchors_out,
  output  fork4_outs_1_valid__anchors_out,
  output  fork4_outs_1_ready__anchors_out,
  output  constant4_outs__data_anchors_out,
  output  constant4_outs_valid__anchors_out,
  output  constant4_outs_ready__anchors_out,
  output [2:0] extsi15_outs__data_anchors_out,
  output  extsi15_outs_valid__anchors_out,
  output  extsi15_outs_ready__anchors_out,
  output [2:0] buffer0_outs__data_anchors_out,
  output  buffer0_outs_valid__anchors_out,
  output  buffer0_outs_ready__anchors_out,
  output [2:0] buffer1_outs__data_anchors_out,
  output  buffer1_outs_valid__anchors_out,
  output  buffer1_outs_ready__anchors_out,
  output [2:0] mux11_outs__data_anchors_out,
  output  mux11_outs_valid__anchors_out,
  output  mux11_outs_ready__anchors_out,
  output [2:0] fork5_outs_0__data_anchors_out,
  output  fork5_outs_0_valid__anchors_out,
  output  fork5_outs_0_ready__anchors_out,
  output [2:0] fork5_outs_1__data_anchors_out,
  output  fork5_outs_1_valid__anchors_out,
  output  fork5_outs_1_ready__anchors_out,
  output [2:0] fork5_outs_2__data_anchors_out,
  output  fork5_outs_2_valid__anchors_out,
  output  fork5_outs_2_ready__anchors_out,
  output [6:0] extsi16_outs__data_anchors_out,
  output  extsi16_outs_valid__anchors_out,
  output  extsi16_outs_ready__anchors_out,
  output [5:0] extsi17_outs__data_anchors_out,
  output  extsi17_outs_valid__anchors_out,
  output  extsi17_outs_ready__anchors_out,
  output [3:0] extsi18_outs__data_anchors_out,
  output  extsi18_outs_valid__anchors_out,
  output  extsi18_outs_ready__anchors_out,
  output [31:0] buffer2_outs__data_anchors_out,
  output  buffer2_outs_valid__anchors_out,
  output  buffer2_outs_ready__anchors_out,
  output [31:0] buffer3_outs__data_anchors_out,
  output  buffer3_outs_valid__anchors_out,
  output  buffer3_outs_ready__anchors_out,
  output [31:0] mux5_outs__data_anchors_out,
  output  mux5_outs_valid__anchors_out,
  output  mux5_outs_ready__anchors_out,
  output [5:0] buffer4_outs__data_anchors_out,
  output  buffer4_outs_valid__anchors_out,
  output  buffer4_outs_ready__anchors_out,
  output [5:0] buffer5_outs__data_anchors_out,
  output  buffer5_outs_valid__anchors_out,
  output  buffer5_outs_ready__anchors_out,
  output [5:0] mux12_outs__data_anchors_out,
  output  mux12_outs_valid__anchors_out,
  output  mux12_outs_ready__anchors_out,
  output [5:0] fork6_outs_0__data_anchors_out,
  output  fork6_outs_0_valid__anchors_out,
  output  fork6_outs_0_ready__anchors_out,
  output [5:0] fork6_outs_1__data_anchors_out,
  output  fork6_outs_1_valid__anchors_out,
  output  fork6_outs_1_ready__anchors_out,
  output [6:0] extsi19_outs__data_anchors_out,
  output  extsi19_outs_valid__anchors_out,
  output  extsi19_outs_ready__anchors_out,
  output [2:0] buffer6_outs__data_anchors_out,
  output  buffer6_outs_valid__anchors_out,
  output  buffer6_outs_ready__anchors_out,
  output [2:0] buffer7_outs__data_anchors_out,
  output  buffer7_outs_valid__anchors_out,
  output  buffer7_outs_ready__anchors_out,
  output [2:0] mux13_outs__data_anchors_out,
  output  mux13_outs_valid__anchors_out,
  output  mux13_outs_ready__anchors_out,
  output [2:0] fork7_outs_0__data_anchors_out,
  output  fork7_outs_0_valid__anchors_out,
  output  fork7_outs_0_ready__anchors_out,
  output [2:0] fork7_outs_1__data_anchors_out,
  output  fork7_outs_1_valid__anchors_out,
  output  fork7_outs_1_ready__anchors_out,
  output [2:0] fork7_outs_2__data_anchors_out,
  output  fork7_outs_2_valid__anchors_out,
  output  fork7_outs_2_ready__anchors_out,
  output [2:0] fork7_outs_3__data_anchors_out,
  output  fork7_outs_3_valid__anchors_out,
  output  fork7_outs_3_ready__anchors_out,
  output [8:0] extsi20_outs__data_anchors_out,
  output  extsi20_outs_valid__anchors_out,
  output  extsi20_outs_ready__anchors_out,
  output [4:0] extsi21_outs__data_anchors_out,
  output  extsi21_outs_valid__anchors_out,
  output  extsi21_outs_ready__anchors_out,
  output [3:0] extsi22_outs__data_anchors_out,
  output  extsi22_outs_valid__anchors_out,
  output  extsi22_outs_ready__anchors_out,
  output  buffer8_outs_valid__anchors_out,
  output  buffer8_outs_ready__anchors_out,
  output  buffer9_outs_valid__anchors_out,
  output  buffer9_outs_ready__anchors_out,
  output  control_merge2_outs_valid__anchors_out,
  output  control_merge2_outs_ready__anchors_out,
  output  control_merge2_index__data_anchors_out,
  output  control_merge2_index_valid__anchors_out,
  output  control_merge2_index_ready__anchors_out,
  output  fork8_outs_0__data_anchors_out,
  output  fork8_outs_0_valid__anchors_out,
  output  fork8_outs_0_ready__anchors_out,
  output  fork8_outs_1__data_anchors_out,
  output  fork8_outs_1_valid__anchors_out,
  output  fork8_outs_1_ready__anchors_out,
  output  fork8_outs_2__data_anchors_out,
  output  fork8_outs_2_valid__anchors_out,
  output  fork8_outs_2_ready__anchors_out,
  output  fork8_outs_3__data_anchors_out,
  output  fork8_outs_3_valid__anchors_out,
  output  fork8_outs_3_ready__anchors_out,
  output  source0_outs_valid__anchors_out,
  output  source0_outs_ready__anchors_out,
  output [5:0] constant5_outs__data_anchors_out,
  output  constant5_outs_valid__anchors_out,
  output  constant5_outs_ready__anchors_out,
  output [8:0] extsi23_outs__data_anchors_out,
  output  extsi23_outs_valid__anchors_out,
  output  extsi23_outs_ready__anchors_out,
  output  source1_outs_valid__anchors_out,
  output  source1_outs_ready__anchors_out,
  output [2:0] constant16_outs__data_anchors_out,
  output  constant16_outs_valid__anchors_out,
  output  constant16_outs_ready__anchors_out,
  output [3:0] extsi24_outs__data_anchors_out,
  output  extsi24_outs_valid__anchors_out,
  output  extsi24_outs_ready__anchors_out,
  output  source2_outs_valid__anchors_out,
  output  source2_outs_ready__anchors_out,
  output [1:0] constant17_outs__data_anchors_out,
  output  constant17_outs_valid__anchors_out,
  output  constant17_outs_ready__anchors_out,
  output [1:0] fork9_outs_0__data_anchors_out,
  output  fork9_outs_0_valid__anchors_out,
  output  fork9_outs_0_ready__anchors_out,
  output [1:0] fork9_outs_1__data_anchors_out,
  output  fork9_outs_1_valid__anchors_out,
  output  fork9_outs_1_ready__anchors_out,
  output [3:0] extui0_outs__data_anchors_out,
  output  extui0_outs_valid__anchors_out,
  output  extui0_outs_ready__anchors_out,
  output [3:0] extsi25_outs__data_anchors_out,
  output  extsi25_outs_valid__anchors_out,
  output  extsi25_outs_ready__anchors_out,
  output [3:0] shli1_result__data_anchors_out,
  output  shli1_result_valid__anchors_out,
  output  shli1_result_ready__anchors_out,
  output [4:0] extsi26_outs__data_anchors_out,
  output  extsi26_outs_valid__anchors_out,
  output  extsi26_outs_ready__anchors_out,
  output [4:0] addi8_result__data_anchors_out,
  output  addi8_result_valid__anchors_out,
  output  addi8_result_ready__anchors_out,
  output [5:0] extsi27_outs__data_anchors_out,
  output  extsi27_outs_valid__anchors_out,
  output  extsi27_outs_ready__anchors_out,
  output [5:0] addi9_result__data_anchors_out,
  output  addi9_result_valid__anchors_out,
  output  addi9_result_ready__anchors_out,
  output [31:0] extsi28_outs__data_anchors_out,
  output  extsi28_outs_valid__anchors_out,
  output  extsi28_outs_ready__anchors_out,
  output [31:0] mc_load0_addrOut__data_anchors_out,
  output  mc_load0_addrOut_valid__anchors_out,
  output  mc_load0_addrOut_ready__anchors_out,
  output [31:0] mc_load0_dataOut__data_anchors_out,
  output  mc_load0_dataOut_valid__anchors_out,
  output  mc_load0_dataOut_ready__anchors_out,
  output [6:0] addi10_result__data_anchors_out,
  output  addi10_result_valid__anchors_out,
  output  addi10_result_ready__anchors_out,
  output [9:0] extsi29_outs__data_anchors_out,
  output  extsi29_outs_valid__anchors_out,
  output  extsi29_outs_ready__anchors_out,
  output [8:0] muli1_result__data_anchors_out,
  output  muli1_result_valid__anchors_out,
  output  muli1_result_ready__anchors_out,
  output [9:0] extsi30_outs__data_anchors_out,
  output  extsi30_outs_valid__anchors_out,
  output  extsi30_outs_ready__anchors_out,
  output [9:0] addi11_result__data_anchors_out,
  output  addi11_result_valid__anchors_out,
  output  addi11_result_ready__anchors_out,
  output [31:0] extsi31_outs__data_anchors_out,
  output  extsi31_outs_valid__anchors_out,
  output  extsi31_outs_ready__anchors_out,
  output [31:0] mc_load1_addrOut__data_anchors_out,
  output  mc_load1_addrOut_valid__anchors_out,
  output  mc_load1_addrOut_ready__anchors_out,
  output [31:0] mc_load1_dataOut__data_anchors_out,
  output  mc_load1_dataOut_valid__anchors_out,
  output  mc_load1_dataOut_ready__anchors_out,
  output [31:0] muli0_result__data_anchors_out,
  output  muli0_result_valid__anchors_out,
  output  muli0_result_ready__anchors_out,
  output [31:0] addi0_result__data_anchors_out,
  output  addi0_result_valid__anchors_out,
  output  addi0_result_ready__anchors_out,
  output [3:0] addi12_result__data_anchors_out,
  output  addi12_result_valid__anchors_out,
  output  addi12_result_ready__anchors_out,
  output [3:0] fork10_outs_0__data_anchors_out,
  output  fork10_outs_0_valid__anchors_out,
  output  fork10_outs_0_ready__anchors_out,
  output [3:0] fork10_outs_1__data_anchors_out,
  output  fork10_outs_1_valid__anchors_out,
  output  fork10_outs_1_ready__anchors_out,
  output [2:0] trunci0_outs__data_anchors_out,
  output  trunci0_outs_valid__anchors_out,
  output  trunci0_outs_ready__anchors_out,
  output  cmpi3_result__data_anchors_out,
  output  cmpi3_result_valid__anchors_out,
  output  cmpi3_result_ready__anchors_out,
  output  fork11_outs_0__data_anchors_out,
  output  fork11_outs_0_valid__anchors_out,
  output  fork11_outs_0_ready__anchors_out,
  output  fork11_outs_1__data_anchors_out,
  output  fork11_outs_1_valid__anchors_out,
  output  fork11_outs_1_ready__anchors_out,
  output  fork11_outs_2__data_anchors_out,
  output  fork11_outs_2_valid__anchors_out,
  output  fork11_outs_2_ready__anchors_out,
  output  fork11_outs_3__data_anchors_out,
  output  fork11_outs_3_valid__anchors_out,
  output  fork11_outs_3_ready__anchors_out,
  output  fork11_outs_4__data_anchors_out,
  output  fork11_outs_4_valid__anchors_out,
  output  fork11_outs_4_ready__anchors_out,
  output [2:0] cond_br0_trueOut__data_anchors_out,
  output  cond_br0_trueOut_valid__anchors_out,
  output  cond_br0_trueOut_ready__anchors_out,
  output [2:0] cond_br0_falseOut__data_anchors_out,
  output  cond_br0_falseOut_valid__anchors_out,
  output  cond_br0_falseOut_ready__anchors_out,
  output [31:0] cond_br4_trueOut__data_anchors_out,
  output  cond_br4_trueOut_valid__anchors_out,
  output  cond_br4_trueOut_ready__anchors_out,
  output [31:0] cond_br4_falseOut__data_anchors_out,
  output  cond_br4_falseOut_valid__anchors_out,
  output  cond_br4_falseOut_ready__anchors_out,
  output [5:0] cond_br1_trueOut__data_anchors_out,
  output  cond_br1_trueOut_valid__anchors_out,
  output  cond_br1_trueOut_ready__anchors_out,
  output [5:0] cond_br1_falseOut__data_anchors_out,
  output  cond_br1_falseOut_valid__anchors_out,
  output  cond_br1_falseOut_ready__anchors_out,
  output [2:0] cond_br2_trueOut__data_anchors_out,
  output  cond_br2_trueOut_valid__anchors_out,
  output  cond_br2_trueOut_ready__anchors_out,
  output [2:0] cond_br2_falseOut__data_anchors_out,
  output  cond_br2_falseOut_valid__anchors_out,
  output  cond_br2_falseOut_ready__anchors_out,
  output  cond_br7_trueOut_valid__anchors_out,
  output  cond_br7_trueOut_ready__anchors_out,
  output  cond_br7_falseOut_valid__anchors_out,
  output  cond_br7_falseOut_ready__anchors_out,
  output [3:0] extsi32_outs__data_anchors_out,
  output  extsi32_outs_valid__anchors_out,
  output  extsi32_outs_ready__anchors_out,
  output  source3_outs_valid__anchors_out,
  output  source3_outs_ready__anchors_out,
  output [2:0] constant18_outs__data_anchors_out,
  output  constant18_outs_valid__anchors_out,
  output  constant18_outs_ready__anchors_out,
  output [3:0] extsi33_outs__data_anchors_out,
  output  extsi33_outs_valid__anchors_out,
  output  extsi33_outs_ready__anchors_out,
  output  source4_outs_valid__anchors_out,
  output  source4_outs_ready__anchors_out,
  output [1:0] constant19_outs__data_anchors_out,
  output  constant19_outs_valid__anchors_out,
  output  constant19_outs_ready__anchors_out,
  output [3:0] extsi34_outs__data_anchors_out,
  output  extsi34_outs_valid__anchors_out,
  output  extsi34_outs_ready__anchors_out,
  output [3:0] addi13_result__data_anchors_out,
  output  addi13_result_valid__anchors_out,
  output  addi13_result_ready__anchors_out,
  output [3:0] fork12_outs_0__data_anchors_out,
  output  fork12_outs_0_valid__anchors_out,
  output  fork12_outs_0_ready__anchors_out,
  output [3:0] fork12_outs_1__data_anchors_out,
  output  fork12_outs_1_valid__anchors_out,
  output  fork12_outs_1_ready__anchors_out,
  output [2:0] trunci1_outs__data_anchors_out,
  output  trunci1_outs_valid__anchors_out,
  output  trunci1_outs_ready__anchors_out,
  output  cmpi4_result__data_anchors_out,
  output  cmpi4_result_valid__anchors_out,
  output  cmpi4_result_ready__anchors_out,
  output  fork13_outs_0__data_anchors_out,
  output  fork13_outs_0_valid__anchors_out,
  output  fork13_outs_0_ready__anchors_out,
  output  fork13_outs_1__data_anchors_out,
  output  fork13_outs_1_valid__anchors_out,
  output  fork13_outs_1_ready__anchors_out,
  output  fork13_outs_2__data_anchors_out,
  output  fork13_outs_2_valid__anchors_out,
  output  fork13_outs_2_ready__anchors_out,
  output  fork13_outs_3__data_anchors_out,
  output  fork13_outs_3_valid__anchors_out,
  output  fork13_outs_3_ready__anchors_out,
  output [2:0] cond_br15_trueOut__data_anchors_out,
  output  cond_br15_trueOut_valid__anchors_out,
  output  cond_br15_trueOut_ready__anchors_out,
  output [2:0] cond_br15_falseOut__data_anchors_out,
  output  cond_br15_falseOut_valid__anchors_out,
  output  cond_br15_falseOut_ready__anchors_out,
  output [31:0] cond_br9_trueOut__data_anchors_out,
  output  cond_br9_trueOut_valid__anchors_out,
  output  cond_br9_trueOut_ready__anchors_out,
  output [31:0] cond_br9_falseOut__data_anchors_out,
  output  cond_br9_falseOut_valid__anchors_out,
  output  cond_br9_falseOut_ready__anchors_out,
  output [5:0] cond_br16_trueOut__data_anchors_out,
  output  cond_br16_trueOut_valid__anchors_out,
  output  cond_br16_trueOut_ready__anchors_out,
  output [5:0] cond_br16_falseOut__data_anchors_out,
  output  cond_br16_falseOut_valid__anchors_out,
  output  cond_br16_falseOut_ready__anchors_out,
  output  cond_br11_trueOut_valid__anchors_out,
  output  cond_br11_trueOut_ready__anchors_out,
  output  cond_br11_falseOut_valid__anchors_out,
  output  cond_br11_falseOut_ready__anchors_out,
  output [1:0] constant20_outs__data_anchors_out,
  output  constant20_outs_valid__anchors_out,
  output  constant20_outs_ready__anchors_out,
  output [31:0] extsi9_outs__data_anchors_out,
  output  extsi9_outs_valid__anchors_out,
  output  extsi9_outs_ready__anchors_out,
  output [5:0] fork14_outs_0__data_anchors_out,
  output  fork14_outs_0_valid__anchors_out,
  output  fork14_outs_0_ready__anchors_out,
  output [5:0] fork14_outs_1__data_anchors_out,
  output  fork14_outs_1_valid__anchors_out,
  output  fork14_outs_1_ready__anchors_out,
  output [6:0] extsi35_outs__data_anchors_out,
  output  extsi35_outs_valid__anchors_out,
  output  extsi35_outs_ready__anchors_out,
  output [31:0] extsi36_outs__data_anchors_out,
  output  extsi36_outs_valid__anchors_out,
  output  extsi36_outs_ready__anchors_out,
  output [31:0] fork15_outs_0__data_anchors_out,
  output  fork15_outs_0_valid__anchors_out,
  output  fork15_outs_0_ready__anchors_out,
  output [31:0] fork15_outs_1__data_anchors_out,
  output  fork15_outs_1_valid__anchors_out,
  output  fork15_outs_1_ready__anchors_out,
  output  fork16_outs_0_valid__anchors_out,
  output  fork16_outs_0_ready__anchors_out,
  output  fork16_outs_1_valid__anchors_out,
  output  fork16_outs_1_ready__anchors_out,
  output  source5_outs_valid__anchors_out,
  output  source5_outs_ready__anchors_out,
  output [5:0] constant21_outs__data_anchors_out,
  output  constant21_outs_valid__anchors_out,
  output  constant21_outs_ready__anchors_out,
  output [6:0] extsi37_outs__data_anchors_out,
  output  extsi37_outs_valid__anchors_out,
  output  extsi37_outs_ready__anchors_out,
  output  source6_outs_valid__anchors_out,
  output  source6_outs_ready__anchors_out,
  output [1:0] constant22_outs__data_anchors_out,
  output  constant22_outs_valid__anchors_out,
  output  constant22_outs_ready__anchors_out,
  output [6:0] extsi38_outs__data_anchors_out,
  output  extsi38_outs_valid__anchors_out,
  output  extsi38_outs_ready__anchors_out,
  output [31:0] mc_store0_addrOut__data_anchors_out,
  output  mc_store0_addrOut_valid__anchors_out,
  output  mc_store0_addrOut_ready__anchors_out,
  output [31:0] mc_store0_dataToMem__data_anchors_out,
  output  mc_store0_dataToMem_valid__anchors_out,
  output  mc_store0_dataToMem_ready__anchors_out,
  output [6:0] addi14_result__data_anchors_out,
  output  addi14_result_valid__anchors_out,
  output  addi14_result_ready__anchors_out,
  output [6:0] fork17_outs_0__data_anchors_out,
  output  fork17_outs_0_valid__anchors_out,
  output  fork17_outs_0_ready__anchors_out,
  output [6:0] fork17_outs_1__data_anchors_out,
  output  fork17_outs_1_valid__anchors_out,
  output  fork17_outs_1_ready__anchors_out,
  output [5:0] trunci2_outs__data_anchors_out,
  output  trunci2_outs_valid__anchors_out,
  output  trunci2_outs_ready__anchors_out,
  output  cmpi5_result__data_anchors_out,
  output  cmpi5_result_valid__anchors_out,
  output  cmpi5_result_ready__anchors_out,
  output  fork18_outs_0__data_anchors_out,
  output  fork18_outs_0_valid__anchors_out,
  output  fork18_outs_0_ready__anchors_out,
  output  fork18_outs_1__data_anchors_out,
  output  fork18_outs_1_valid__anchors_out,
  output  fork18_outs_1_ready__anchors_out,
  output  fork18_outs_2__data_anchors_out,
  output  fork18_outs_2_valid__anchors_out,
  output  fork18_outs_2_ready__anchors_out,
  output [5:0] cond_br17_trueOut__data_anchors_out,
  output  cond_br17_trueOut_valid__anchors_out,
  output  cond_br17_trueOut_ready__anchors_out,
  output [5:0] cond_br17_falseOut__data_anchors_out,
  output  cond_br17_falseOut_valid__anchors_out,
  output  cond_br17_falseOut_ready__anchors_out,
  output  cond_br13_trueOut_valid__anchors_out,
  output  cond_br13_trueOut_ready__anchors_out,
  output  cond_br13_falseOut_valid__anchors_out,
  output  cond_br13_falseOut_ready__anchors_out,
  output [31:0] cond_br14_trueOut__data_anchors_out,
  output  cond_br14_trueOut_valid__anchors_out,
  output  cond_br14_trueOut_ready__anchors_out,
  output [31:0] cond_br14_falseOut__data_anchors_out,
  output  cond_br14_falseOut_valid__anchors_out,
  output  cond_br14_falseOut_ready__anchors_out,
  output  fork19_outs_0_valid__anchors_out,
  output  fork19_outs_0_ready__anchors_out,
  output  fork19_outs_1_valid__anchors_out,
  output  fork19_outs_1_ready__anchors_out,
  output  fork19_outs_2_valid__anchors_out,
  output  fork19_outs_2_ready__anchors_out
);
  wire  mem_controller0_loadEn;
  wire [31:0] mem_controller0_loadAddr;
  wire  mem_controller0_storeEn;
  wire [31:0] mem_controller0_storeAddr;
  wire [31:0] mem_controller0_storeData;
  wire  mem_controller1_loadEn;
  wire [31:0] mem_controller1_loadAddr;
  wire  mem_controller1_storeEn;
  wire [31:0] mem_controller1_storeAddr;
  wire [31:0] mem_controller1_storeData;
  wire  mem_controller2_loadEn;
  wire [31:0] mem_controller2_loadAddr;
  wire  mem_controller2_storeEn;
  wire [31:0] mem_controller2_storeAddr;
  wire [31:0] mem_controller2_storeData;

  // module outputs
  assign out0 = cond_br14_falseOut__data_anchors_out;
  assign out0_valid = cond_br14_falseOut_valid__anchors_out;
  assign cond_br14_falseOut_ready = out0_ready;
  assign orig_end_valid = mem_controller2_memEnd_valid__anchors_out;
  assign mem_controller2_memEnd_ready = orig_end_ready;
  assign filter_end_valid = mem_controller1_memEnd_valid__anchors_out;
  assign mem_controller1_memEnd_ready = filter_end_ready;
  assign sol_end_valid = mem_controller0_memEnd_valid__anchors_out;
  assign mem_controller0_memEnd_ready = sol_end_ready;
  assign end_valid = fork0_outs_1_valid__anchors_out;
  assign fork0_outs_1_ready = end_ready;
  assign orig_loadEn = mem_controller2_loadEn;
  assign orig_loadAddr = mem_controller2_loadAddr;
  assign orig_storeEn = mem_controller2_storeEn;
  assign orig_storeAddr = mem_controller2_storeAddr;
  assign orig_storeData = mem_controller2_storeData;
  assign filter_loadEn = mem_controller1_loadEn;
  assign filter_loadAddr = mem_controller1_loadAddr;
  assign filter_storeEn = mem_controller1_storeEn;
  assign filter_storeAddr = mem_controller1_storeAddr;
  assign filter_storeData = mem_controller1_storeData;
  assign sol_loadEn = mem_controller0_loadEn;
  assign sol_loadAddr = mem_controller0_loadAddr;
  assign sol_storeEn = mem_controller0_storeEn;
  assign sol_storeAddr = mem_controller0_storeAddr;
  assign sol_storeData = mem_controller0_storeData;


fork_dataless #(.SIZE(3)) fork0(
.clk (clk),
.ins_ready (start_ready),
.ins_valid (start_valid),
.outs_ready ({fork0_outs_2_ready__anchors_in, fork0_outs_1_ready__anchors_in, fork0_outs_0_ready__anchors_in}),
.outs_valid ({fork0_outs_2_valid__anchors_out, fork0_outs_1_valid__anchors_out, fork0_outs_0_valid__anchors_out}),
.rst (rst)
);

mem_controller_loadless #(.NUM_CONTROLS(1), .NUM_STORES(1), .DATA_TYPE(32), .ADDR_TYPE(32)) mem_controller0(
.clk (clk),
.ctrl ({extsi9_outs__data_anchors_in}),
.ctrlEnd_ready (fork19_outs_0_ready__anchors_out),
.ctrlEnd_valid (fork19_outs_0_valid__anchors_in),
.ctrl_ready ({extsi9_outs_ready__anchors_out}),
.ctrl_valid ({extsi9_outs_valid__anchors_in}),
.loadAddr (mem_controller0_loadAddr),
.loadData (sol_loadData),
.loadEn (mem_controller0_loadEn),
.memEnd_ready (mem_controller0_memEnd_ready),
.memEnd_valid (mem_controller0_memEnd_valid),
.memStart_ready (sol_start_ready),
.memStart_valid (sol_start_valid),
.rst (rst),
.stAddr ({mc_store0_addrOut}),
.stAddr_ready ({mc_store0_addrOut_ready}),
.stAddr_valid ({mc_store0_addrOut_valid}),
.stData ({mc_store0_dataToMem}),
.stData_ready ({mc_store0_dataToMem_ready}),
.stData_valid ({mc_store0_dataToMem_valid}),
.storeAddr (mem_controller0_storeAddr),
.storeData (mem_controller0_storeData),
.storeEn (mem_controller0_storeEn)
);

mem_controller_storeless #(.NUM_LOADS(1), .DATA_TYPE(32), .ADDR_TYPE(32)) mem_controller1(
.clk (clk),
.ctrlEnd_ready (fork19_outs_1_ready__anchors_out),
.ctrlEnd_valid (fork19_outs_1_valid__anchors_in),
.ldAddr ({mc_load0_addrOut}),
.ldAddr_ready ({mc_load0_addrOut_ready}),
.ldAddr_valid ({mc_load0_addrOut_valid}),
.ldData ({mem_controller1_ldData_0}),
.ldData_ready ({mem_controller1_ldData_0_ready}),
.ldData_valid ({mem_controller1_ldData_0_valid}),
.loadAddr (mem_controller1_loadAddr),
.loadData (filter_loadData),
.loadEn (mem_controller1_loadEn),
.memEnd_ready (mem_controller1_memEnd_ready),
.memEnd_valid (mem_controller1_memEnd_valid),
.memStart_ready (filter_start_ready),
.memStart_valid (filter_start_valid),
.rst (rst),
.storeAddr (mem_controller1_storeAddr),
.storeData (mem_controller1_storeData),
.storeEn (mem_controller1_storeEn)
);

mem_controller_storeless #(.NUM_LOADS(1), .DATA_TYPE(32), .ADDR_TYPE(32)) mem_controller2(
.clk (clk),
.ctrlEnd_ready (fork19_outs_2_ready__anchors_out),
.ctrlEnd_valid (fork19_outs_2_valid__anchors_in),
.ldAddr ({mc_load1_addrOut}),
.ldAddr_ready ({mc_load1_addrOut_ready}),
.ldAddr_valid ({mc_load1_addrOut_valid}),
.ldData ({mem_controller2_ldData_0}),
.ldData_ready ({mem_controller2_ldData_0_ready}),
.ldData_valid ({mem_controller2_ldData_0_valid}),
.loadAddr (mem_controller2_loadAddr),
.loadData (orig_loadData),
.loadEn (mem_controller2_loadEn),
.memEnd_ready (mem_controller2_memEnd_ready),
.memEnd_valid (mem_controller2_memEnd_valid),
.memStart_ready (orig_start_ready),
.memStart_valid (orig_start_valid),
.rst (rst),
.storeAddr (mem_controller2_storeAddr),
.storeData (mem_controller2_storeData),
.storeEn (mem_controller2_storeEn)
);

handshake_constant_0 #(.DATA_WIDTH(1)) constant1(
.clk (clk),
.ctrl_ready (fork0_outs_0_ready__anchors_out),
.ctrl_valid (fork0_outs_0_valid__anchors_in),
.outs (constant1_outs__data_anchors_out),
.outs_ready (constant1_outs_ready__anchors_in),
.outs_valid (constant1_outs_valid__anchors_out),
.rst (rst)
);

extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(6)) extsi12(
.clk (clk),
.ins (constant1_outs__data_anchors_in),
.ins_ready (constant1_outs_ready__anchors_out),
.ins_valid (constant1_outs_valid__anchors_in),
.outs (extsi12_outs__data_anchors_out),
.outs_ready (extsi12_outs_ready__anchors_in),
.outs_valid (extsi12_outs_valid__anchors_out),
.rst (rst)
);

oehb #(.DATA_TYPE(6)) buffer18(
.clk (clk),
.ins (cond_br17_trueOut__data_anchors_in),
.ins_ready (cond_br17_trueOut_ready__anchors_out),
.ins_valid (cond_br17_trueOut_valid__anchors_in),
.outs (buffer18_outs__data_anchors_out),
.outs_ready (buffer18_outs_ready__anchors_in),
.outs_valid (buffer18_outs_valid__anchors_out),
.rst (rst)
);

tehb #(.DATA_TYPE(6)) buffer19(
.clk (clk),
.ins (buffer18_outs__data_anchors_in),
.ins_ready (buffer18_outs_ready__anchors_out),
.ins_valid (buffer18_outs_valid__anchors_in),
.outs (buffer19_outs__data_anchors_out),
.outs_ready (buffer19_outs_ready__anchors_in),
.outs_valid (buffer19_outs_valid__anchors_out),
.rst (rst)
);

mux #(.SIZE(2), .DATA_TYPE(6), .SELECT_TYPE(1)) mux8(
.clk (clk),
.index (control_merge0_index),
.index_ready (control_merge0_index_ready__anchors_out),
.index_valid (control_merge0_index_valid),
.ins ({buffer19_outs__data_anchors_in, extsi12_outs__data_anchors_in}),
.ins_ready ({buffer19_outs_ready__anchors_out, extsi12_outs_ready__anchors_out}),
.ins_valid ({buffer19_outs_valid__anchors_in, extsi12_outs_valid__anchors_in}),
.outs (mux8_outs__data_anchors_out),
.outs_ready (mux8_outs_ready__anchors_in),
.outs_valid (mux8_outs_valid__anchors_out),
.rst (rst)
);

oehb_dataless buffer20(
.clk (clk),
.ins_ready (cond_br13_trueOut_ready__anchors_out),
.ins_valid (cond_br13_trueOut_valid__anchors_in),
.outs_ready (buffer20_outs_ready__anchors_in),
.outs_valid (buffer20_outs_valid__anchors_out),
.rst (rst)
);

tehb_dataless buffer21(
.clk (clk),
.ins_ready (buffer20_outs_ready__anchors_out),
.ins_valid (buffer20_outs_valid__anchors_in),
.outs_ready (buffer21_outs_ready__anchors_in),
.outs_valid (buffer21_outs_valid__anchors_out),
.rst (rst)
);

control_merge_dataless #(.SIZE(2), .INDEX_TYPE(1)) control_merge0(
.clk (clk),
.index (control_merge0_index),
.index_ready (control_merge0_index_ready__anchors_in),
.index_valid (control_merge0_index_valid),
.ins_ready ({buffer21_outs_ready__anchors_out, fork0_outs_2_ready__anchors_out}),
.ins_valid ({buffer21_outs_valid__anchors_in, fork0_outs_2_valid__anchors_in}),
.outs_ready (control_merge0_outs_ready__anchors_in),
.outs_valid (control_merge0_outs_valid__anchors_out),
.rst (rst)
);

fork_dataless #(.SIZE(2)) fork1(
.clk (clk),
.ins_ready (control_merge0_outs_ready__anchors_out),
.ins_valid (control_merge0_outs_valid__anchors_in),
.outs_ready ({fork1_outs_1_ready__anchors_in, fork1_outs_0_ready__anchors_in}),
.outs_valid ({fork1_outs_1_valid__anchors_out, fork1_outs_0_valid__anchors_out}),
.rst (rst)
);

handshake_constant_0 #(.DATA_WIDTH(1)) constant3(
.clk (clk),
.ctrl_ready (fork1_outs_0_ready__anchors_out),
.ctrl_valid (fork1_outs_0_valid__anchors_in),
.outs (constant3_outs__data_anchors_out),
.outs_ready (constant3_outs_ready__anchors_in),
.outs_valid (constant3_outs_valid__anchors_out),
.rst (rst)
);

fork_type #(.SIZE(2), .DATA_TYPE(1)) fork2(
.clk (clk),
.ins (constant3_outs__data_anchors_in),
.ins_ready (constant3_outs_ready__anchors_out),
.ins_valid (constant3_outs_valid__anchors_in),
.outs ({fork2_outs_1__data_anchors_out, fork2_outs_0__data_anchors_out}),
.outs_ready ({fork2_outs_1_ready__anchors_in, fork2_outs_0_ready__anchors_in}),
.outs_valid ({fork2_outs_1_valid__anchors_out, fork2_outs_0_valid__anchors_out}),
.rst (rst)
);

extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(3)) extsi13(
.clk (clk),
.ins (fork2_outs_0__data_anchors_in),
.ins_ready (fork2_outs_0_ready__anchors_out),
.ins_valid (fork2_outs_0_valid__anchors_in),
.outs (extsi13_outs__data_anchors_out),
.outs_ready (extsi13_outs_ready__anchors_in),
.outs_valid (extsi13_outs_valid__anchors_out),
.rst (rst)
);

extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(32)) extsi14(
.clk (clk),
.ins (fork2_outs_1__data_anchors_in),
.ins_ready (fork2_outs_1_ready__anchors_out),
.ins_valid (fork2_outs_1_valid__anchors_in),
.outs (extsi14_outs__data_anchors_out),
.outs_ready (extsi14_outs_ready__anchors_in),
.outs_valid (extsi14_outs_valid__anchors_out),
.rst (rst)
);

oehb #(.DATA_TYPE(3)) buffer10(
.clk (clk),
.ins (cond_br15_trueOut__data_anchors_in),
.ins_ready (cond_br15_trueOut_ready__anchors_out),
.ins_valid (cond_br15_trueOut_valid__anchors_in),
.outs (buffer10_outs__data_anchors_out),
.outs_ready (buffer10_outs_ready__anchors_in),
.outs_valid (buffer10_outs_valid__anchors_out),
.rst (rst)
);

tehb #(.DATA_TYPE(3)) buffer11(
.clk (clk),
.ins (buffer10_outs__data_anchors_in),
.ins_ready (buffer10_outs_ready__anchors_out),
.ins_valid (buffer10_outs_valid__anchors_in),
.outs (buffer11_outs__data_anchors_out),
.outs_ready (buffer11_outs_ready__anchors_in),
.outs_valid (buffer11_outs_valid__anchors_out),
.rst (rst)
);

mux #(.SIZE(2), .DATA_TYPE(3), .SELECT_TYPE(1)) mux9(
.clk (clk),
.index (fork3_outs_1__data_anchors_in),
.index_ready (fork3_outs_1_ready__anchors_out),
.index_valid (fork3_outs_1_valid__anchors_in),
.ins ({buffer11_outs__data_anchors_in, extsi13_outs__data_anchors_in}),
.ins_ready ({buffer11_outs_ready__anchors_out, extsi13_outs_ready__anchors_out}),
.ins_valid ({buffer11_outs_valid__anchors_in, extsi13_outs_valid__anchors_in}),
.outs (mux9_outs__data_anchors_out),
.outs_ready (mux9_outs_ready__anchors_in),
.outs_valid (mux9_outs_valid__anchors_out),
.rst (rst)
);

oehb #(.DATA_TYPE(32)) buffer12(
.clk (clk),
.ins (cond_br9_trueOut__data_anchors_in),
.ins_ready (cond_br9_trueOut_ready__anchors_out),
.ins_valid (cond_br9_trueOut_valid__anchors_in),
.outs (buffer12_outs__data_anchors_out),
.outs_ready (buffer12_outs_ready__anchors_in),
.outs_valid (buffer12_outs_valid__anchors_out),
.rst (rst)
);

tehb #(.DATA_TYPE(32)) buffer13(
.clk (clk),
.ins (buffer12_outs__data_anchors_in),
.ins_ready (buffer12_outs_ready__anchors_out),
.ins_valid (buffer12_outs_valid__anchors_in),
.outs (buffer13_outs__data_anchors_out),
.outs_ready (buffer13_outs_ready__anchors_in),
.outs_valid (buffer13_outs_valid__anchors_out),
.rst (rst)
);

mux #(.SIZE(2), .DATA_TYPE(32), .SELECT_TYPE(1)) mux2(
.clk (clk),
.index (fork3_outs_2__data_anchors_in),
.index_ready (fork3_outs_2_ready__anchors_out),
.index_valid (fork3_outs_2_valid__anchors_in),
.ins ({buffer13_outs__data_anchors_in, extsi14_outs__data_anchors_in}),
.ins_ready ({buffer13_outs_ready__anchors_out, extsi14_outs_ready__anchors_out}),
.ins_valid ({buffer13_outs_valid__anchors_in, extsi14_outs_valid__anchors_in}),
.outs (mux2_outs__data_anchors_out),
.outs_ready (mux2_outs_ready__anchors_in),
.outs_valid (mux2_outs_valid__anchors_out),
.rst (rst)
);

oehb #(.DATA_TYPE(6)) buffer14(
.clk (clk),
.ins (cond_br16_trueOut__data_anchors_in),
.ins_ready (cond_br16_trueOut_ready__anchors_out),
.ins_valid (cond_br16_trueOut_valid__anchors_in),
.outs (buffer14_outs__data_anchors_out),
.outs_ready (buffer14_outs_ready__anchors_in),
.outs_valid (buffer14_outs_valid__anchors_out),
.rst (rst)
);

tehb #(.DATA_TYPE(6)) buffer15(
.clk (clk),
.ins (buffer14_outs__data_anchors_in),
.ins_ready (buffer14_outs_ready__anchors_out),
.ins_valid (buffer14_outs_valid__anchors_in),
.outs (buffer15_outs__data_anchors_out),
.outs_ready (buffer15_outs_ready__anchors_in),
.outs_valid (buffer15_outs_valid__anchors_out),
.rst (rst)
);

mux #(.SIZE(2), .DATA_TYPE(6), .SELECT_TYPE(1)) mux10(
.clk (clk),
.index (fork3_outs_0__data_anchors_in),
.index_ready (fork3_outs_0_ready__anchors_out),
.index_valid (fork3_outs_0_valid__anchors_in),
.ins ({buffer15_outs__data_anchors_in, mux8_outs__data_anchors_in}),
.ins_ready ({buffer15_outs_ready__anchors_out, mux8_outs_ready__anchors_out}),
.ins_valid ({buffer15_outs_valid__anchors_in, mux8_outs_valid__anchors_in}),
.outs (mux10_outs__data_anchors_out),
.outs_ready (mux10_outs_ready__anchors_in),
.outs_valid (mux10_outs_valid__anchors_out),
.rst (rst)
);

oehb_dataless buffer16(
.clk (clk),
.ins_ready (cond_br11_trueOut_ready__anchors_out),
.ins_valid (cond_br11_trueOut_valid__anchors_in),
.outs_ready (buffer16_outs_ready__anchors_in),
.outs_valid (buffer16_outs_valid__anchors_out),
.rst (rst)
);

tehb_dataless buffer17(
.clk (clk),
.ins_ready (buffer16_outs_ready__anchors_out),
.ins_valid (buffer16_outs_valid__anchors_in),
.outs_ready (buffer17_outs_ready__anchors_in),
.outs_valid (buffer17_outs_valid__anchors_out),
.rst (rst)
);

control_merge_dataless #(.SIZE(2), .INDEX_TYPE(1)) control_merge1(
.clk (clk),
.index (control_merge1_index),
.index_ready (control_merge1_index_ready__anchors_in),
.index_valid (control_merge1_index_valid),
.ins_ready ({buffer17_outs_ready__anchors_out, fork1_outs_1_ready__anchors_out}),
.ins_valid ({buffer17_outs_valid__anchors_in, fork1_outs_1_valid__anchors_in}),
.outs_ready (control_merge1_outs_ready__anchors_in),
.outs_valid (control_merge1_outs_valid__anchors_out),
.rst (rst)
);

fork_type #(.SIZE(3), .DATA_TYPE(1)) fork3(
.clk (clk),
.ins (control_merge1_index__data_anchors_in),
.ins_ready (control_merge1_index_ready__anchors_out),
.ins_valid (control_merge1_index_valid__anchors_in),
.outs ({fork3_outs_2__data_anchors_out, fork3_outs_1__data_anchors_out, fork3_outs_0__data_anchors_out}),
.outs_ready ({fork3_outs_2_ready__anchors_in, fork3_outs_1_ready__anchors_in, fork3_outs_0_ready__anchors_in}),
.outs_valid ({fork3_outs_2_valid__anchors_out, fork3_outs_1_valid__anchors_out, fork3_outs_0_valid__anchors_out}),
.rst (rst)
);

fork_dataless #(.SIZE(2)) fork4(
.clk (clk),
.ins_ready (control_merge1_outs_ready__anchors_out),
.ins_valid (control_merge1_outs_valid__anchors_in),
.outs_ready ({fork4_outs_1_ready__anchors_in, fork4_outs_0_ready__anchors_in}),
.outs_valid ({fork4_outs_1_valid__anchors_out, fork4_outs_0_valid__anchors_out}),
.rst (rst)
);

handshake_constant_0 #(.DATA_WIDTH(1)) constant4(
.clk (clk),
.ctrl_ready (fork4_outs_0_ready__anchors_out),
.ctrl_valid (fork4_outs_0_valid__anchors_in),
.outs (constant4_outs__data_anchors_out),
.outs_ready (constant4_outs_ready__anchors_in),
.outs_valid (constant4_outs_valid__anchors_out),
.rst (rst)
);

extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(3)) extsi15(
.clk (clk),
.ins (constant4_outs__data_anchors_in),
.ins_ready (constant4_outs_ready__anchors_out),
.ins_valid (constant4_outs_valid__anchors_in),
.outs (extsi15_outs__data_anchors_out),
.outs_ready (extsi15_outs_ready__anchors_in),
.outs_valid (extsi15_outs_valid__anchors_out),
.rst (rst)
);

oehb #(.DATA_TYPE(3)) buffer0(
.clk (clk),
.ins (cond_br0_trueOut__data_anchors_in),
.ins_ready (cond_br0_trueOut_ready__anchors_out),
.ins_valid (cond_br0_trueOut_valid__anchors_in),
.outs (buffer0_outs__data_anchors_out),
.outs_ready (buffer0_outs_ready__anchors_in),
.outs_valid (buffer0_outs_valid__anchors_out),
.rst (rst)
);

tehb #(.DATA_TYPE(3)) buffer1(
.clk (clk),
.ins (buffer0_outs__data_anchors_in),
.ins_ready (buffer0_outs_ready__anchors_out),
.ins_valid (buffer0_outs_valid__anchors_in),
.outs (buffer1_outs__data_anchors_out),
.outs_ready (buffer1_outs_ready__anchors_in),
.outs_valid (buffer1_outs_valid__anchors_out),
.rst (rst)
);

mux #(.SIZE(2), .DATA_TYPE(3), .SELECT_TYPE(1)) mux11(
.clk (clk),
.index (fork8_outs_2__data_anchors_in),
.index_ready (fork8_outs_2_ready__anchors_out),
.index_valid (fork8_outs_2_valid__anchors_in),
.ins ({buffer1_outs__data_anchors_in, extsi15_outs__data_anchors_in}),
.ins_ready ({buffer1_outs_ready__anchors_out, extsi15_outs_ready__anchors_out}),
.ins_valid ({buffer1_outs_valid__anchors_in, extsi15_outs_valid__anchors_in}),
.outs (mux11_outs__data_anchors_out),
.outs_ready (mux11_outs_ready__anchors_in),
.outs_valid (mux11_outs_valid__anchors_out),
.rst (rst)
);

fork_type #(.SIZE(3), .DATA_TYPE(3)) fork5(
.clk (clk),
.ins (mux11_outs__data_anchors_in),
.ins_ready (mux11_outs_ready__anchors_out),
.ins_valid (mux11_outs_valid__anchors_in),
.outs ({fork5_outs_2__data_anchors_out, fork5_outs_1__data_anchors_out, fork5_outs_0__data_anchors_out}),
.outs_ready ({fork5_outs_2_ready__anchors_in, fork5_outs_1_ready__anchors_in, fork5_outs_0_ready__anchors_in}),
.outs_valid ({fork5_outs_2_valid__anchors_out, fork5_outs_1_valid__anchors_out, fork5_outs_0_valid__anchors_out}),
.rst (rst)
);

extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(7)) extsi16(
.clk (clk),
.ins (fork5_outs_0__data_anchors_in),
.ins_ready (fork5_outs_0_ready__anchors_out),
.ins_valid (fork5_outs_0_valid__anchors_in),
.outs (extsi16_outs__data_anchors_out),
.outs_ready (extsi16_outs_ready__anchors_in),
.outs_valid (extsi16_outs_valid__anchors_out),
.rst (rst)
);

extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(6)) extsi17(
.clk (clk),
.ins (fork5_outs_1__data_anchors_in),
.ins_ready (fork5_outs_1_ready__anchors_out),
.ins_valid (fork5_outs_1_valid__anchors_in),
.outs (extsi17_outs__data_anchors_out),
.outs_ready (extsi17_outs_ready__anchors_in),
.outs_valid (extsi17_outs_valid__anchors_out),
.rst (rst)
);

extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(4)) extsi18(
.clk (clk),
.ins (fork5_outs_2__data_anchors_in),
.ins_ready (fork5_outs_2_ready__anchors_out),
.ins_valid (fork5_outs_2_valid__anchors_in),
.outs (extsi18_outs__data_anchors_out),
.outs_ready (extsi18_outs_ready__anchors_in),
.outs_valid (extsi18_outs_valid__anchors_out),
.rst (rst)
);

oehb #(.DATA_TYPE(32)) buffer2(
.clk (clk),
.ins (cond_br4_trueOut__data_anchors_in),
.ins_ready (cond_br4_trueOut_ready__anchors_out),
.ins_valid (cond_br4_trueOut_valid__anchors_in),
.outs (buffer2_outs__data_anchors_out),
.outs_ready (buffer2_outs_ready__anchors_in),
.outs_valid (buffer2_outs_valid__anchors_out),
.rst (rst)
);

tehb #(.DATA_TYPE(32)) buffer3(
.clk (clk),
.ins (buffer2_outs__data_anchors_in),
.ins_ready (buffer2_outs_ready__anchors_out),
.ins_valid (buffer2_outs_valid__anchors_in),
.outs (buffer3_outs__data_anchors_out),
.outs_ready (buffer3_outs_ready__anchors_in),
.outs_valid (buffer3_outs_valid__anchors_out),
.rst (rst)
);

mux #(.SIZE(2), .DATA_TYPE(32), .SELECT_TYPE(1)) mux5(
.clk (clk),
.index (fork8_outs_3__data_anchors_in),
.index_ready (fork8_outs_3_ready__anchors_out),
.index_valid (fork8_outs_3_valid__anchors_in),
.ins ({buffer3_outs__data_anchors_in, mux2_outs__data_anchors_in}),
.ins_ready ({buffer3_outs_ready__anchors_out, mux2_outs_ready__anchors_out}),
.ins_valid ({buffer3_outs_valid__anchors_in, mux2_outs_valid__anchors_in}),
.outs (mux5_outs__data_anchors_out),
.outs_ready (mux5_outs_ready__anchors_in),
.outs_valid (mux5_outs_valid__anchors_out),
.rst (rst)
);

oehb #(.DATA_TYPE(6)) buffer4(
.clk (clk),
.ins (cond_br1_trueOut__data_anchors_in),
.ins_ready (cond_br1_trueOut_ready__anchors_out),
.ins_valid (cond_br1_trueOut_valid__anchors_in),
.outs (buffer4_outs__data_anchors_out),
.outs_ready (buffer4_outs_ready__anchors_in),
.outs_valid (buffer4_outs_valid__anchors_out),
.rst (rst)
);

tehb #(.DATA_TYPE(6)) buffer5(
.clk (clk),
.ins (buffer4_outs__data_anchors_in),
.ins_ready (buffer4_outs_ready__anchors_out),
.ins_valid (buffer4_outs_valid__anchors_in),
.outs (buffer5_outs__data_anchors_out),
.outs_ready (buffer5_outs_ready__anchors_in),
.outs_valid (buffer5_outs_valid__anchors_out),
.rst (rst)
);

mux #(.SIZE(2), .DATA_TYPE(6), .SELECT_TYPE(1)) mux12(
.clk (clk),
.index (fork8_outs_0__data_anchors_in),
.index_ready (fork8_outs_0_ready__anchors_out),
.index_valid (fork8_outs_0_valid__anchors_in),
.ins ({buffer5_outs__data_anchors_in, mux10_outs__data_anchors_in}),
.ins_ready ({buffer5_outs_ready__anchors_out, mux10_outs_ready__anchors_out}),
.ins_valid ({buffer5_outs_valid__anchors_in, mux10_outs_valid__anchors_in}),
.outs (mux12_outs__data_anchors_out),
.outs_ready (mux12_outs_ready__anchors_in),
.outs_valid (mux12_outs_valid__anchors_out),
.rst (rst)
);

fork_type #(.SIZE(2), .DATA_TYPE(6)) fork6(
.clk (clk),
.ins (mux12_outs__data_anchors_in),
.ins_ready (mux12_outs_ready__anchors_out),
.ins_valid (mux12_outs_valid__anchors_in),
.outs ({fork6_outs_1__data_anchors_out, fork6_outs_0__data_anchors_out}),
.outs_ready ({fork6_outs_1_ready__anchors_in, fork6_outs_0_ready__anchors_in}),
.outs_valid ({fork6_outs_1_valid__anchors_out, fork6_outs_0_valid__anchors_out}),
.rst (rst)
);

extsi #(.INPUT_TYPE(6), .OUTPUT_TYPE(7)) extsi19(
.clk (clk),
.ins (fork6_outs_1__data_anchors_in),
.ins_ready (fork6_outs_1_ready__anchors_out),
.ins_valid (fork6_outs_1_valid__anchors_in),
.outs (extsi19_outs__data_anchors_out),
.outs_ready (extsi19_outs_ready__anchors_in),
.outs_valid (extsi19_outs_valid__anchors_out),
.rst (rst)
);

oehb #(.DATA_TYPE(3)) buffer6(
.clk (clk),
.ins (cond_br2_trueOut__data_anchors_in),
.ins_ready (cond_br2_trueOut_ready__anchors_out),
.ins_valid (cond_br2_trueOut_valid__anchors_in),
.outs (buffer6_outs__data_anchors_out),
.outs_ready (buffer6_outs_ready__anchors_in),
.outs_valid (buffer6_outs_valid__anchors_out),
.rst (rst)
);

tehb #(.DATA_TYPE(3)) buffer7(
.clk (clk),
.ins (buffer6_outs__data_anchors_in),
.ins_ready (buffer6_outs_ready__anchors_out),
.ins_valid (buffer6_outs_valid__anchors_in),
.outs (buffer7_outs__data_anchors_out),
.outs_ready (buffer7_outs_ready__anchors_in),
.outs_valid (buffer7_outs_valid__anchors_out),
.rst (rst)
);

mux #(.SIZE(2), .DATA_TYPE(3), .SELECT_TYPE(1)) mux13(
.clk (clk),
.index (fork8_outs_1__data_anchors_in),
.index_ready (fork8_outs_1_ready__anchors_out),
.index_valid (fork8_outs_1_valid__anchors_in),
.ins ({buffer7_outs__data_anchors_in, mux9_outs__data_anchors_in}),
.ins_ready ({buffer7_outs_ready__anchors_out, mux9_outs_ready__anchors_out}),
.ins_valid ({buffer7_outs_valid__anchors_in, mux9_outs_valid__anchors_in}),
.outs (mux13_outs__data_anchors_out),
.outs_ready (mux13_outs_ready__anchors_in),
.outs_valid (mux13_outs_valid__anchors_out),
.rst (rst)
);

fork_type #(.SIZE(4), .DATA_TYPE(3)) fork7(
.clk (clk),
.ins (mux13_outs__data_anchors_in),
.ins_ready (mux13_outs_ready__anchors_out),
.ins_valid (mux13_outs_valid__anchors_in),
.outs ({fork7_outs_3__data_anchors_out, fork7_outs_2__data_anchors_out, fork7_outs_1__data_anchors_out, fork7_outs_0__data_anchors_out}),
.outs_ready ({fork7_outs_3_ready__anchors_in, fork7_outs_2_ready__anchors_in, fork7_outs_1_ready__anchors_in, fork7_outs_0_ready__anchors_in}),
.outs_valid ({fork7_outs_3_valid__anchors_out, fork7_outs_2_valid__anchors_out, fork7_outs_1_valid__anchors_out, fork7_outs_0_valid__anchors_out}),
.rst (rst)
);

extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(9)) extsi20(
.clk (clk),
.ins (fork7_outs_1__data_anchors_in),
.ins_ready (fork7_outs_1_ready__anchors_out),
.ins_valid (fork7_outs_1_valid__anchors_in),
.outs (extsi20_outs__data_anchors_out),
.outs_ready (extsi20_outs_ready__anchors_in),
.outs_valid (extsi20_outs_valid__anchors_out),
.rst (rst)
);

extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(5)) extsi21(
.clk (clk),
.ins (fork7_outs_2__data_anchors_in),
.ins_ready (fork7_outs_2_ready__anchors_out),
.ins_valid (fork7_outs_2_valid__anchors_in),
.outs (extsi21_outs__data_anchors_out),
.outs_ready (extsi21_outs_ready__anchors_in),
.outs_valid (extsi21_outs_valid__anchors_out),
.rst (rst)
);

extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(4)) extsi22(
.clk (clk),
.ins (fork7_outs_3__data_anchors_in),
.ins_ready (fork7_outs_3_ready__anchors_out),
.ins_valid (fork7_outs_3_valid__anchors_in),
.outs (extsi22_outs__data_anchors_out),
.outs_ready (extsi22_outs_ready__anchors_in),
.outs_valid (extsi22_outs_valid__anchors_out),
.rst (rst)
);

oehb_dataless buffer8(
.clk (clk),
.ins_ready (cond_br7_trueOut_ready__anchors_out),
.ins_valid (cond_br7_trueOut_valid__anchors_in),
.outs_ready (buffer8_outs_ready__anchors_in),
.outs_valid (buffer8_outs_valid__anchors_out),
.rst (rst)
);

tehb_dataless buffer9(
.clk (clk),
.ins_ready (buffer8_outs_ready__anchors_out),
.ins_valid (buffer8_outs_valid__anchors_in),
.outs_ready (buffer9_outs_ready__anchors_in),
.outs_valid (buffer9_outs_valid__anchors_out),
.rst (rst)
);

control_merge_dataless #(.SIZE(2), .INDEX_TYPE(1)) control_merge2(
.clk (clk),
.index (control_merge2_index),
.index_ready (control_merge2_index_ready__anchors_in),
.index_valid (control_merge2_index_valid),
.ins_ready ({buffer9_outs_ready__anchors_out, fork4_outs_1_ready__anchors_out}),
.ins_valid ({buffer9_outs_valid__anchors_in, fork4_outs_1_valid__anchors_in}),
.outs_ready (control_merge2_outs_ready__anchors_in),
.outs_valid (control_merge2_outs_valid__anchors_out),
.rst (rst)
);

fork_type #(.SIZE(4), .DATA_TYPE(1)) fork8(
.clk (clk),
.ins (control_merge2_index__data_anchors_in),
.ins_ready (control_merge2_index_ready__anchors_out),
.ins_valid (control_merge2_index_valid__anchors_in),
.outs ({fork8_outs_3__data_anchors_out, fork8_outs_2__data_anchors_out, fork8_outs_1__data_anchors_out, fork8_outs_0__data_anchors_out}),
.outs_ready ({fork8_outs_3_ready__anchors_in, fork8_outs_2_ready__anchors_in, fork8_outs_1_ready__anchors_in, fork8_outs_0_ready__anchors_in}),
.outs_valid ({fork8_outs_3_valid__anchors_out, fork8_outs_2_valid__anchors_out, fork8_outs_1_valid__anchors_out, fork8_outs_0_valid__anchors_out}),
.rst (rst)
);

source source0(
.clk (clk),
.outs_ready (source0_outs_ready__anchors_in),
.outs_valid (source0_outs_valid__anchors_out),
.rst (rst)
);

handshake_constant_1 #(.DATA_WIDTH(6)) constant5(
.clk (clk),
.ctrl_ready (source0_outs_ready__anchors_out),
.ctrl_valid (source0_outs_valid__anchors_in),
.outs (constant5_outs__data_anchors_out),
.outs_ready (constant5_outs_ready__anchors_in),
.outs_valid (constant5_outs_valid__anchors_out),
.rst (rst)
);

extsi #(.INPUT_TYPE(6), .OUTPUT_TYPE(9)) extsi23(
.clk (clk),
.ins (constant5_outs__data_anchors_in),
.ins_ready (constant5_outs_ready__anchors_out),
.ins_valid (constant5_outs_valid__anchors_in),
.outs (extsi23_outs__data_anchors_out),
.outs_ready (extsi23_outs_ready__anchors_in),
.outs_valid (extsi23_outs_valid__anchors_out),
.rst (rst)
);

source source1(
.clk (clk),
.outs_ready (source1_outs_ready__anchors_in),
.outs_valid (source1_outs_valid__anchors_out),
.rst (rst)
);

handshake_constant_2 #(.DATA_WIDTH(3)) constant16(
.clk (clk),
.ctrl_ready (source1_outs_ready__anchors_out),
.ctrl_valid (source1_outs_valid__anchors_in),
.outs (constant16_outs__data_anchors_out),
.outs_ready (constant16_outs_ready__anchors_in),
.outs_valid (constant16_outs_valid__anchors_out),
.rst (rst)
);

extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(4)) extsi24(
.clk (clk),
.ins (constant16_outs__data_anchors_in),
.ins_ready (constant16_outs_ready__anchors_out),
.ins_valid (constant16_outs_valid__anchors_in),
.outs (extsi24_outs__data_anchors_out),
.outs_ready (extsi24_outs_ready__anchors_in),
.outs_valid (extsi24_outs_valid__anchors_out),
.rst (rst)
);

source source2(
.clk (clk),
.outs_ready (source2_outs_ready__anchors_in),
.outs_valid (source2_outs_valid__anchors_out),
.rst (rst)
);

handshake_constant_3 #(.DATA_WIDTH(2)) constant17(
.clk (clk),
.ctrl_ready (source2_outs_ready__anchors_out),
.ctrl_valid (source2_outs_valid__anchors_in),
.outs (constant17_outs__data_anchors_out),
.outs_ready (constant17_outs_ready__anchors_in),
.outs_valid (constant17_outs_valid__anchors_out),
.rst (rst)
);

fork_type #(.SIZE(2), .DATA_TYPE(2)) fork9(
.clk (clk),
.ins (constant17_outs__data_anchors_in),
.ins_ready (constant17_outs_ready__anchors_out),
.ins_valid (constant17_outs_valid__anchors_in),
.outs ({fork9_outs_1__data_anchors_out, fork9_outs_0__data_anchors_out}),
.outs_ready ({fork9_outs_1_ready__anchors_in, fork9_outs_0_ready__anchors_in}),
.outs_valid ({fork9_outs_1_valid__anchors_out, fork9_outs_0_valid__anchors_out}),
.rst (rst)
);

extui #(.INPUT_TYPE(2), .OUTPUT_TYPE(4)) extui0(
.clk (clk),
.ins (fork9_outs_0__data_anchors_in),
.ins_ready (fork9_outs_0_ready__anchors_out),
.ins_valid (fork9_outs_0_valid__anchors_in),
.outs (extui0_outs__data_anchors_out),
.outs_ready (extui0_outs_ready__anchors_in),
.outs_valid (extui0_outs_valid__anchors_out),
.rst (rst)
);

extsi #(.INPUT_TYPE(2), .OUTPUT_TYPE(4)) extsi25(
.clk (clk),
.ins (fork9_outs_1__data_anchors_in),
.ins_ready (fork9_outs_1_ready__anchors_out),
.ins_valid (fork9_outs_1_valid__anchors_in),
.outs (extsi25_outs__data_anchors_out),
.outs_ready (extsi25_outs_ready__anchors_in),
.outs_valid (extsi25_outs_valid__anchors_out),
.rst (rst)
);

shli #(.DATA_TYPE(4)) shli1(
.clk (clk),
.lhs (extsi22_outs__data_anchors_in),
.lhs_ready (extsi22_outs_ready__anchors_out),
.lhs_valid (extsi22_outs_valid__anchors_in),
.result (shli1_result__data_anchors_out),
.result_ready (shli1_result_ready__anchors_in),
.result_valid (shli1_result_valid__anchors_out),
.rhs (extui0_outs__data_anchors_in),
.rhs_ready (extui0_outs_ready__anchors_out),
.rhs_valid (extui0_outs_valid__anchors_in),
.rst (rst)
);

extsi #(.INPUT_TYPE(4), .OUTPUT_TYPE(5)) extsi26(
.clk (clk),
.ins (shli1_result__data_anchors_in),
.ins_ready (shli1_result_ready__anchors_out),
.ins_valid (shli1_result_valid__anchors_in),
.outs (extsi26_outs__data_anchors_out),
.outs_ready (extsi26_outs_ready__anchors_in),
.outs_valid (extsi26_outs_valid__anchors_out),
.rst (rst)
);

addi #(.DATA_TYPE(5)) addi8(
.clk (clk),
.lhs (extsi21_outs__data_anchors_in),
.lhs_ready (extsi21_outs_ready__anchors_out),
.lhs_valid (extsi21_outs_valid__anchors_in),
.result (addi8_result__data_anchors_out),
.result_ready (addi8_result_ready__anchors_in),
.result_valid (addi8_result_valid__anchors_out),
.rhs (extsi26_outs__data_anchors_in),
.rhs_ready (extsi26_outs_ready__anchors_out),
.rhs_valid (extsi26_outs_valid__anchors_in),
.rst (rst)
);

extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(6)) extsi27(
.clk (clk),
.ins (addi8_result__data_anchors_in),
.ins_ready (addi8_result_ready__anchors_out),
.ins_valid (addi8_result_valid__anchors_in),
.outs (extsi27_outs__data_anchors_out),
.outs_ready (extsi27_outs_ready__anchors_in),
.outs_valid (extsi27_outs_valid__anchors_out),
.rst (rst)
);

addi #(.DATA_TYPE(6)) addi9(
.clk (clk),
.lhs (extsi17_outs__data_anchors_in),
.lhs_ready (extsi17_outs_ready__anchors_out),
.lhs_valid (extsi17_outs_valid__anchors_in),
.result (addi9_result__data_anchors_out),
.result_ready (addi9_result_ready__anchors_in),
.result_valid (addi9_result_valid__anchors_out),
.rhs (extsi27_outs__data_anchors_in),
.rhs_ready (extsi27_outs_ready__anchors_out),
.rhs_valid (extsi27_outs_valid__anchors_in),
.rst (rst)
);

extsi #(.INPUT_TYPE(6), .OUTPUT_TYPE(32)) extsi28(
.clk (clk),
.ins (addi9_result__data_anchors_in),
.ins_ready (addi9_result_ready__anchors_out),
.ins_valid (addi9_result_valid__anchors_in),
.outs (extsi28_outs__data_anchors_out),
.outs_ready (extsi28_outs_ready__anchors_in),
.outs_valid (extsi28_outs_valid__anchors_out),
.rst (rst)
);

mc_load #(.DATA_TYPE(32), .ADDR_TYPE(32)) mc_load0(
.addrIn (extsi28_outs__data_anchors_in),
.addrIn_ready (extsi28_outs_ready__anchors_out),
.addrIn_valid (extsi28_outs_valid__anchors_in),
.addrOut (mc_load0_addrOut),
.addrOut_ready (mc_load0_addrOut_ready),
.addrOut_valid (mc_load0_addrOut_valid),
.clk (clk),
.dataFromMem (mem_controller1_ldData_0__data_anchors_in),
.dataFromMem_ready (mem_controller1_ldData_0_ready__anchors_out),
.dataFromMem_valid (mem_controller1_ldData_0_valid__anchors_in),
.dataOut (mc_load0_dataOut),
.dataOut_ready (mc_load0_dataOut_ready),
.dataOut_valid (mc_load0_dataOut_valid),
.rst (rst)
);

addi #(.DATA_TYPE(7)) addi10(
.clk (clk),
.lhs (extsi16_outs__data_anchors_in),
.lhs_ready (extsi16_outs_ready__anchors_out),
.lhs_valid (extsi16_outs_valid__anchors_in),
.result (addi10_result__data_anchors_out),
.result_ready (addi10_result_ready__anchors_in),
.result_valid (addi10_result_valid__anchors_out),
.rhs (extsi19_outs__data_anchors_in),
.rhs_ready (extsi19_outs_ready__anchors_out),
.rhs_valid (extsi19_outs_valid__anchors_in),
.rst (rst)
);

extsi #(.INPUT_TYPE(7), .OUTPUT_TYPE(10)) extsi29(
.clk (clk),
.ins (addi10_result__data_anchors_in),
.ins_ready (addi10_result_ready__anchors_out),
.ins_valid (addi10_result_valid__anchors_in),
.outs (extsi29_outs__data_anchors_out),
.outs_ready (extsi29_outs_ready__anchors_in),
.outs_valid (extsi29_outs_valid__anchors_out),
.rst (rst)
);

muli #(.DATA_TYPE(9)) muli1(
.clk (clk),
.lhs (extsi20_outs__data_anchors_in),
.lhs_ready (extsi20_outs_ready__anchors_out),
.lhs_valid (extsi20_outs_valid__anchors_in),
.result (muli1_result__data_anchors_out),
.result_ready (muli1_result_ready__anchors_in),
.result_valid (muli1_result_valid__anchors_out),
.rhs (extsi23_outs__data_anchors_in),
.rhs_ready (extsi23_outs_ready__anchors_out),
.rhs_valid (extsi23_outs_valid__anchors_in),
.rst (rst)
);

extsi #(.INPUT_TYPE(9), .OUTPUT_TYPE(10)) extsi30(
.clk (clk),
.ins (muli1_result__data_anchors_in),
.ins_ready (muli1_result_ready__anchors_out),
.ins_valid (muli1_result_valid__anchors_in),
.outs (extsi30_outs__data_anchors_out),
.outs_ready (extsi30_outs_ready__anchors_in),
.outs_valid (extsi30_outs_valid__anchors_out),
.rst (rst)
);

addi #(.DATA_TYPE(10)) addi11(
.clk (clk),
.lhs (extsi29_outs__data_anchors_in),
.lhs_ready (extsi29_outs_ready__anchors_out),
.lhs_valid (extsi29_outs_valid__anchors_in),
.result (addi11_result__data_anchors_out),
.result_ready (addi11_result_ready__anchors_in),
.result_valid (addi11_result_valid__anchors_out),
.rhs (extsi30_outs__data_anchors_in),
.rhs_ready (extsi30_outs_ready__anchors_out),
.rhs_valid (extsi30_outs_valid__anchors_in),
.rst (rst)
);

extsi #(.INPUT_TYPE(10), .OUTPUT_TYPE(32)) extsi31(
.clk (clk),
.ins (addi11_result__data_anchors_in),
.ins_ready (addi11_result_ready__anchors_out),
.ins_valid (addi11_result_valid__anchors_in),
.outs (extsi31_outs__data_anchors_out),
.outs_ready (extsi31_outs_ready__anchors_in),
.outs_valid (extsi31_outs_valid__anchors_out),
.rst (rst)
);

mc_load #(.DATA_TYPE(32), .ADDR_TYPE(32)) mc_load1(
.addrIn (extsi31_outs__data_anchors_in),
.addrIn_ready (extsi31_outs_ready__anchors_out),
.addrIn_valid (extsi31_outs_valid__anchors_in),
.addrOut (mc_load1_addrOut),
.addrOut_ready (mc_load1_addrOut_ready),
.addrOut_valid (mc_load1_addrOut_valid),
.clk (clk),
.dataFromMem (mem_controller2_ldData_0__data_anchors_in),
.dataFromMem_ready (mem_controller2_ldData_0_ready__anchors_out),
.dataFromMem_valid (mem_controller2_ldData_0_valid__anchors_in),
.dataOut (mc_load1_dataOut),
.dataOut_ready (mc_load1_dataOut_ready),
.dataOut_valid (mc_load1_dataOut_valid),
.rst (rst)
);

muli #(.DATA_TYPE(32)) muli0(
.clk (clk),
.lhs (mc_load0_dataOut),
.lhs_ready (mc_load0_dataOut_ready),
.lhs_valid (mc_load0_dataOut_valid),
.result (muli0_result__data_anchors_out),
.result_ready (muli0_result_ready__anchors_in),
.result_valid (muli0_result_valid__anchors_out),
.rhs (mc_load1_dataOut),
.rhs_ready (mc_load1_dataOut_ready),
.rhs_valid (mc_load1_dataOut_valid),
.rst (rst)
);

addi #(.DATA_TYPE(32)) addi0(
.clk (clk),
.lhs (mux5_outs__data_anchors_in),
.lhs_ready (mux5_outs_ready__anchors_out),
.lhs_valid (mux5_outs_valid__anchors_in),
.result (addi0_result__data_anchors_out),
.result_ready (addi0_result_ready__anchors_in),
.result_valid (addi0_result_valid__anchors_out),
.rhs (muli0_result__data_anchors_in),
.rhs_ready (muli0_result_ready__anchors_out),
.rhs_valid (muli0_result_valid__anchors_in),
.rst (rst)
);

addi #(.DATA_TYPE(4)) addi12(
.clk (clk),
.lhs (extsi18_outs__data_anchors_in),
.lhs_ready (extsi18_outs_ready__anchors_out),
.lhs_valid (extsi18_outs_valid__anchors_in),
.result (addi12_result__data_anchors_out),
.result_ready (addi12_result_ready__anchors_in),
.result_valid (addi12_result_valid__anchors_out),
.rhs (extsi25_outs__data_anchors_in),
.rhs_ready (extsi25_outs_ready__anchors_out),
.rhs_valid (extsi25_outs_valid__anchors_in),
.rst (rst)
);

fork_type #(.SIZE(2), .DATA_TYPE(4)) fork10(
.clk (clk),
.ins (addi12_result__data_anchors_in),
.ins_ready (addi12_result_ready__anchors_out),
.ins_valid (addi12_result_valid__anchors_in),
.outs ({fork10_outs_1__data_anchors_out, fork10_outs_0__data_anchors_out}),
.outs_ready ({fork10_outs_1_ready__anchors_in, fork10_outs_0_ready__anchors_in}),
.outs_valid ({fork10_outs_1_valid__anchors_out, fork10_outs_0_valid__anchors_out}),
.rst (rst)
);

trunci #(.INPUT_TYPE(4), .OUTPUT_TYPE(3)) trunci0(
.clk (clk),
.ins (fork10_outs_0__data_anchors_in),
.ins_ready (fork10_outs_0_ready__anchors_out),
.ins_valid (fork10_outs_0_valid__anchors_in),
.outs (trunci0_outs__data_anchors_out),
.outs_ready (trunci0_outs_ready__anchors_in),
.outs_valid (trunci0_outs_valid__anchors_out),
.rst (rst)
);

handshake_cmpi_0 #(.DATA_TYPE(4)) cmpi3(
.clk (clk),
.lhs (fork10_outs_1__data_anchors_in),
.lhs_ready (fork10_outs_1_ready__anchors_out),
.lhs_valid (fork10_outs_1_valid__anchors_in),
.result (cmpi3_result__data_anchors_out),
.result_ready (cmpi3_result_ready__anchors_in),
.result_valid (cmpi3_result_valid__anchors_out),
.rhs (extsi24_outs__data_anchors_in),
.rhs_ready (extsi24_outs_ready__anchors_out),
.rhs_valid (extsi24_outs_valid__anchors_in),
.rst (rst)
);

fork_type #(.SIZE(5), .DATA_TYPE(1)) fork11(
.clk (clk),
.ins (cmpi3_result__data_anchors_in),
.ins_ready (cmpi3_result_ready__anchors_out),
.ins_valid (cmpi3_result_valid__anchors_in),
.outs ({fork11_outs_4__data_anchors_out, fork11_outs_3__data_anchors_out, fork11_outs_2__data_anchors_out, fork11_outs_1__data_anchors_out, fork11_outs_0__data_anchors_out}),
.outs_ready ({fork11_outs_4_ready__anchors_in, fork11_outs_3_ready__anchors_in, fork11_outs_2_ready__anchors_in, fork11_outs_1_ready__anchors_in, fork11_outs_0_ready__anchors_in}),
.outs_valid ({fork11_outs_4_valid__anchors_out, fork11_outs_3_valid__anchors_out, fork11_outs_2_valid__anchors_out, fork11_outs_1_valid__anchors_out, fork11_outs_0_valid__anchors_out}),
.rst (rst)
);

cond_br #(.DATA_TYPE(3)) cond_br0(
.clk (clk),
.condition (fork11_outs_0__data_anchors_in),
.condition_ready (fork11_outs_0_ready__anchors_out),
.condition_valid (fork11_outs_0_valid__anchors_in),
.data (trunci0_outs__data_anchors_in),
.data_ready (trunci0_outs_ready__anchors_out),
.data_valid (trunci0_outs_valid__anchors_in),
.falseOut (cond_br0_falseOut__data_anchors_out),
.falseOut_ready (cond_br0_falseOut_ready__anchors_in),
.falseOut_valid (cond_br0_falseOut_valid__anchors_out),
.rst (rst),
.trueOut (cond_br0_trueOut__data_anchors_out),
.trueOut_ready (cond_br0_trueOut_ready__anchors_in),
.trueOut_valid (cond_br0_trueOut_valid__anchors_out)
);

sink #(.DATA_TYPE(3)) sink0(
.clk (clk),
.ins (cond_br0_falseOut__data_anchors_in),
.ins_ready (cond_br0_falseOut_ready__anchors_out),
.ins_valid (cond_br0_falseOut_valid__anchors_in),
.rst (rst)
);

cond_br #(.DATA_TYPE(32)) cond_br4(
.clk (clk),
.condition (fork11_outs_3__data_anchors_in),
.condition_ready (fork11_outs_3_ready__anchors_out),
.condition_valid (fork11_outs_3_valid__anchors_in),
.data (addi0_result__data_anchors_in),
.data_ready (addi0_result_ready__anchors_out),
.data_valid (addi0_result_valid__anchors_in),
.falseOut (cond_br4_falseOut__data_anchors_out),
.falseOut_ready (cond_br4_falseOut_ready__anchors_in),
.falseOut_valid (cond_br4_falseOut_valid__anchors_out),
.rst (rst),
.trueOut (cond_br4_trueOut__data_anchors_out),
.trueOut_ready (cond_br4_trueOut_ready__anchors_in),
.trueOut_valid (cond_br4_trueOut_valid__anchors_out)
);

cond_br #(.DATA_TYPE(6)) cond_br1(
.clk (clk),
.condition (fork11_outs_1__data_anchors_in),
.condition_ready (fork11_outs_1_ready__anchors_out),
.condition_valid (fork11_outs_1_valid__anchors_in),
.data (fork6_outs_0__data_anchors_in),
.data_ready (fork6_outs_0_ready__anchors_out),
.data_valid (fork6_outs_0_valid__anchors_in),
.falseOut (cond_br1_falseOut__data_anchors_out),
.falseOut_ready (cond_br1_falseOut_ready__anchors_in),
.falseOut_valid (cond_br1_falseOut_valid__anchors_out),
.rst (rst),
.trueOut (cond_br1_trueOut__data_anchors_out),
.trueOut_ready (cond_br1_trueOut_ready__anchors_in),
.trueOut_valid (cond_br1_trueOut_valid__anchors_out)
);

cond_br #(.DATA_TYPE(3)) cond_br2(
.clk (clk),
.condition (fork11_outs_2__data_anchors_in),
.condition_ready (fork11_outs_2_ready__anchors_out),
.condition_valid (fork11_outs_2_valid__anchors_in),
.data (fork7_outs_0__data_anchors_in),
.data_ready (fork7_outs_0_ready__anchors_out),
.data_valid (fork7_outs_0_valid__anchors_in),
.falseOut (cond_br2_falseOut__data_anchors_out),
.falseOut_ready (cond_br2_falseOut_ready__anchors_in),
.falseOut_valid (cond_br2_falseOut_valid__anchors_out),
.rst (rst),
.trueOut (cond_br2_trueOut__data_anchors_out),
.trueOut_ready (cond_br2_trueOut_ready__anchors_in),
.trueOut_valid (cond_br2_trueOut_valid__anchors_out)
);

cond_br_dataless cond_br7(
.clk (clk),
.condition (fork11_outs_4__data_anchors_in),
.condition_ready (fork11_outs_4_ready__anchors_out),
.condition_valid (fork11_outs_4_valid__anchors_in),
.data_ready (control_merge2_outs_ready__anchors_out),
.data_valid (control_merge2_outs_valid__anchors_in),
.falseOut_ready (cond_br7_falseOut_ready__anchors_in),
.falseOut_valid (cond_br7_falseOut_valid__anchors_out),
.rst (rst),
.trueOut_ready (cond_br7_trueOut_ready__anchors_in),
.trueOut_valid (cond_br7_trueOut_valid__anchors_out)
);

extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(4)) extsi32(
.clk (clk),
.ins (cond_br2_falseOut__data_anchors_in),
.ins_ready (cond_br2_falseOut_ready__anchors_out),
.ins_valid (cond_br2_falseOut_valid__anchors_in),
.outs (extsi32_outs__data_anchors_out),
.outs_ready (extsi32_outs_ready__anchors_in),
.outs_valid (extsi32_outs_valid__anchors_out),
.rst (rst)
);

source source3(
.clk (clk),
.outs_ready (source3_outs_ready__anchors_in),
.outs_valid (source3_outs_valid__anchors_out),
.rst (rst)
);

handshake_constant_2 #(.DATA_WIDTH(3)) constant18(
.clk (clk),
.ctrl_ready (source3_outs_ready__anchors_out),
.ctrl_valid (source3_outs_valid__anchors_in),
.outs (constant18_outs__data_anchors_out),
.outs_ready (constant18_outs_ready__anchors_in),
.outs_valid (constant18_outs_valid__anchors_out),
.rst (rst)
);

extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(4)) extsi33(
.clk (clk),
.ins (constant18_outs__data_anchors_in),
.ins_ready (constant18_outs_ready__anchors_out),
.ins_valid (constant18_outs_valid__anchors_in),
.outs (extsi33_outs__data_anchors_out),
.outs_ready (extsi33_outs_ready__anchors_in),
.outs_valid (extsi33_outs_valid__anchors_out),
.rst (rst)
);

source source4(
.clk (clk),
.outs_ready (source4_outs_ready__anchors_in),
.outs_valid (source4_outs_valid__anchors_out),
.rst (rst)
);

handshake_constant_3 #(.DATA_WIDTH(2)) constant19(
.clk (clk),
.ctrl_ready (source4_outs_ready__anchors_out),
.ctrl_valid (source4_outs_valid__anchors_in),
.outs (constant19_outs__data_anchors_out),
.outs_ready (constant19_outs_ready__anchors_in),
.outs_valid (constant19_outs_valid__anchors_out),
.rst (rst)
);

extsi #(.INPUT_TYPE(2), .OUTPUT_TYPE(4)) extsi34(
.clk (clk),
.ins (constant19_outs__data_anchors_in),
.ins_ready (constant19_outs_ready__anchors_out),
.ins_valid (constant19_outs_valid__anchors_in),
.outs (extsi34_outs__data_anchors_out),
.outs_ready (extsi34_outs_ready__anchors_in),
.outs_valid (extsi34_outs_valid__anchors_out),
.rst (rst)
);

addi #(.DATA_TYPE(4)) addi13(
.clk (clk),
.lhs (extsi32_outs__data_anchors_in),
.lhs_ready (extsi32_outs_ready__anchors_out),
.lhs_valid (extsi32_outs_valid__anchors_in),
.result (addi13_result__data_anchors_out),
.result_ready (addi13_result_ready__anchors_in),
.result_valid (addi13_result_valid__anchors_out),
.rhs (extsi34_outs__data_anchors_in),
.rhs_ready (extsi34_outs_ready__anchors_out),
.rhs_valid (extsi34_outs_valid__anchors_in),
.rst (rst)
);

fork_type #(.SIZE(2), .DATA_TYPE(4)) fork12(
.clk (clk),
.ins (addi13_result__data_anchors_in),
.ins_ready (addi13_result_ready__anchors_out),
.ins_valid (addi13_result_valid__anchors_in),
.outs ({fork12_outs_1__data_anchors_out, fork12_outs_0__data_anchors_out}),
.outs_ready ({fork12_outs_1_ready__anchors_in, fork12_outs_0_ready__anchors_in}),
.outs_valid ({fork12_outs_1_valid__anchors_out, fork12_outs_0_valid__anchors_out}),
.rst (rst)
);

trunci #(.INPUT_TYPE(4), .OUTPUT_TYPE(3)) trunci1(
.clk (clk),
.ins (fork12_outs_0__data_anchors_in),
.ins_ready (fork12_outs_0_ready__anchors_out),
.ins_valid (fork12_outs_0_valid__anchors_in),
.outs (trunci1_outs__data_anchors_out),
.outs_ready (trunci1_outs_ready__anchors_in),
.outs_valid (trunci1_outs_valid__anchors_out),
.rst (rst)
);

handshake_cmpi_0 #(.DATA_TYPE(4)) cmpi4(
.clk (clk),
.lhs (fork12_outs_1__data_anchors_in),
.lhs_ready (fork12_outs_1_ready__anchors_out),
.lhs_valid (fork12_outs_1_valid__anchors_in),
.result (cmpi4_result__data_anchors_out),
.result_ready (cmpi4_result_ready__anchors_in),
.result_valid (cmpi4_result_valid__anchors_out),
.rhs (extsi33_outs__data_anchors_in),
.rhs_ready (extsi33_outs_ready__anchors_out),
.rhs_valid (extsi33_outs_valid__anchors_in),
.rst (rst)
);

fork_type #(.SIZE(4), .DATA_TYPE(1)) fork13(
.clk (clk),
.ins (cmpi4_result__data_anchors_in),
.ins_ready (cmpi4_result_ready__anchors_out),
.ins_valid (cmpi4_result_valid__anchors_in),
.outs ({fork13_outs_3__data_anchors_out, fork13_outs_2__data_anchors_out, fork13_outs_1__data_anchors_out, fork13_outs_0__data_anchors_out}),
.outs_ready ({fork13_outs_3_ready__anchors_in, fork13_outs_2_ready__anchors_in, fork13_outs_1_ready__anchors_in, fork13_outs_0_ready__anchors_in}),
.outs_valid ({fork13_outs_3_valid__anchors_out, fork13_outs_2_valid__anchors_out, fork13_outs_1_valid__anchors_out, fork13_outs_0_valid__anchors_out}),
.rst (rst)
);

cond_br #(.DATA_TYPE(3)) cond_br15(
.clk (clk),
.condition (fork13_outs_0__data_anchors_in),
.condition_ready (fork13_outs_0_ready__anchors_out),
.condition_valid (fork13_outs_0_valid__anchors_in),
.data (trunci1_outs__data_anchors_in),
.data_ready (trunci1_outs_ready__anchors_out),
.data_valid (trunci1_outs_valid__anchors_in),
.falseOut (cond_br15_falseOut__data_anchors_out),
.falseOut_ready (cond_br15_falseOut_ready__anchors_in),
.falseOut_valid (cond_br15_falseOut_valid__anchors_out),
.rst (rst),
.trueOut (cond_br15_trueOut__data_anchors_out),
.trueOut_ready (cond_br15_trueOut_ready__anchors_in),
.trueOut_valid (cond_br15_trueOut_valid__anchors_out)
);

sink #(.DATA_TYPE(3)) sink2(
.clk (clk),
.ins (cond_br15_falseOut__data_anchors_in),
.ins_ready (cond_br15_falseOut_ready__anchors_out),
.ins_valid (cond_br15_falseOut_valid__anchors_in),
.rst (rst)
);

cond_br #(.DATA_TYPE(32)) cond_br9(
.clk (clk),
.condition (fork13_outs_2__data_anchors_in),
.condition_ready (fork13_outs_2_ready__anchors_out),
.condition_valid (fork13_outs_2_valid__anchors_in),
.data (cond_br4_falseOut__data_anchors_in),
.data_ready (cond_br4_falseOut_ready__anchors_out),
.data_valid (cond_br4_falseOut_valid__anchors_in),
.falseOut (cond_br9_falseOut__data_anchors_out),
.falseOut_ready (cond_br9_falseOut_ready__anchors_in),
.falseOut_valid (cond_br9_falseOut_valid__anchors_out),
.rst (rst),
.trueOut (cond_br9_trueOut__data_anchors_out),
.trueOut_ready (cond_br9_trueOut_ready__anchors_in),
.trueOut_valid (cond_br9_trueOut_valid__anchors_out)
);

cond_br #(.DATA_TYPE(6)) cond_br16(
.clk (clk),
.condition (fork13_outs_1__data_anchors_in),
.condition_ready (fork13_outs_1_ready__anchors_out),
.condition_valid (fork13_outs_1_valid__anchors_in),
.data (cond_br1_falseOut__data_anchors_in),
.data_ready (cond_br1_falseOut_ready__anchors_out),
.data_valid (cond_br1_falseOut_valid__anchors_in),
.falseOut (cond_br16_falseOut__data_anchors_out),
.falseOut_ready (cond_br16_falseOut_ready__anchors_in),
.falseOut_valid (cond_br16_falseOut_valid__anchors_out),
.rst (rst),
.trueOut (cond_br16_trueOut__data_anchors_out),
.trueOut_ready (cond_br16_trueOut_ready__anchors_in),
.trueOut_valid (cond_br16_trueOut_valid__anchors_out)
);

cond_br_dataless cond_br11(
.clk (clk),
.condition (fork13_outs_3__data_anchors_in),
.condition_ready (fork13_outs_3_ready__anchors_out),
.condition_valid (fork13_outs_3_valid__anchors_in),
.data_ready (cond_br7_falseOut_ready__anchors_out),
.data_valid (cond_br7_falseOut_valid__anchors_in),
.falseOut_ready (cond_br11_falseOut_ready__anchors_in),
.falseOut_valid (cond_br11_falseOut_valid__anchors_out),
.rst (rst),
.trueOut_ready (cond_br11_trueOut_ready__anchors_in),
.trueOut_valid (cond_br11_trueOut_valid__anchors_out)
);

handshake_constant_3 #(.DATA_WIDTH(2)) constant20(
.clk (clk),
.ctrl_ready (fork16_outs_0_ready__anchors_out),
.ctrl_valid (fork16_outs_0_valid__anchors_in),
.outs (constant20_outs__data_anchors_out),
.outs_ready (constant20_outs_ready__anchors_in),
.outs_valid (constant20_outs_valid__anchors_out),
.rst (rst)
);

extsi #(.INPUT_TYPE(2), .OUTPUT_TYPE(32)) extsi9(
.clk (clk),
.ins (constant20_outs__data_anchors_in),
.ins_ready (constant20_outs_ready__anchors_out),
.ins_valid (constant20_outs_valid__anchors_in),
.outs (extsi9_outs__data_anchors_out),
.outs_ready (extsi9_outs_ready__anchors_in),
.outs_valid (extsi9_outs_valid__anchors_out),
.rst (rst)
);

fork_type #(.SIZE(2), .DATA_TYPE(6)) fork14(
.clk (clk),
.ins (cond_br16_falseOut__data_anchors_in),
.ins_ready (cond_br16_falseOut_ready__anchors_out),
.ins_valid (cond_br16_falseOut_valid__anchors_in),
.outs ({fork14_outs_1__data_anchors_out, fork14_outs_0__data_anchors_out}),
.outs_ready ({fork14_outs_1_ready__anchors_in, fork14_outs_0_ready__anchors_in}),
.outs_valid ({fork14_outs_1_valid__anchors_out, fork14_outs_0_valid__anchors_out}),
.rst (rst)
);

extsi #(.INPUT_TYPE(6), .OUTPUT_TYPE(7)) extsi35(
.clk (clk),
.ins (fork14_outs_0__data_anchors_in),
.ins_ready (fork14_outs_0_ready__anchors_out),
.ins_valid (fork14_outs_0_valid__anchors_in),
.outs (extsi35_outs__data_anchors_out),
.outs_ready (extsi35_outs_ready__anchors_in),
.outs_valid (extsi35_outs_valid__anchors_out),
.rst (rst)
);

extsi #(.INPUT_TYPE(6), .OUTPUT_TYPE(32)) extsi36(
.clk (clk),
.ins (fork14_outs_1__data_anchors_in),
.ins_ready (fork14_outs_1_ready__anchors_out),
.ins_valid (fork14_outs_1_valid__anchors_in),
.outs (extsi36_outs__data_anchors_out),
.outs_ready (extsi36_outs_ready__anchors_in),
.outs_valid (extsi36_outs_valid__anchors_out),
.rst (rst)
);

fork_type #(.SIZE(2), .DATA_TYPE(32)) fork15(
.clk (clk),
.ins (cond_br9_falseOut__data_anchors_in),
.ins_ready (cond_br9_falseOut_ready__anchors_out),
.ins_valid (cond_br9_falseOut_valid__anchors_in),
.outs ({fork15_outs_1__data_anchors_out, fork15_outs_0__data_anchors_out}),
.outs_ready ({fork15_outs_1_ready__anchors_in, fork15_outs_0_ready__anchors_in}),
.outs_valid ({fork15_outs_1_valid__anchors_out, fork15_outs_0_valid__anchors_out}),
.rst (rst)
);

fork_dataless #(.SIZE(2)) fork16(
.clk (clk),
.ins_ready (cond_br11_falseOut_ready__anchors_out),
.ins_valid (cond_br11_falseOut_valid__anchors_in),
.outs_ready ({fork16_outs_1_ready__anchors_in, fork16_outs_0_ready__anchors_in}),
.outs_valid ({fork16_outs_1_valid__anchors_out, fork16_outs_0_valid__anchors_out}),
.rst (rst)
);

source source5(
.clk (clk),
.outs_ready (source5_outs_ready__anchors_in),
.outs_valid (source5_outs_valid__anchors_out),
.rst (rst)
);

handshake_constant_4 #(.DATA_WIDTH(6)) constant21(
.clk (clk),
.ctrl_ready (source5_outs_ready__anchors_out),
.ctrl_valid (source5_outs_valid__anchors_in),
.outs (constant21_outs__data_anchors_out),
.outs_ready (constant21_outs_ready__anchors_in),
.outs_valid (constant21_outs_valid__anchors_out),
.rst (rst)
);

extsi #(.INPUT_TYPE(6), .OUTPUT_TYPE(7)) extsi37(
.clk (clk),
.ins (constant21_outs__data_anchors_in),
.ins_ready (constant21_outs_ready__anchors_out),
.ins_valid (constant21_outs_valid__anchors_in),
.outs (extsi37_outs__data_anchors_out),
.outs_ready (extsi37_outs_ready__anchors_in),
.outs_valid (extsi37_outs_valid__anchors_out),
.rst (rst)
);

source source6(
.clk (clk),
.outs_ready (source6_outs_ready__anchors_in),
.outs_valid (source6_outs_valid__anchors_out),
.rst (rst)
);

handshake_constant_3 #(.DATA_WIDTH(2)) constant22(
.clk (clk),
.ctrl_ready (source6_outs_ready__anchors_out),
.ctrl_valid (source6_outs_valid__anchors_in),
.outs (constant22_outs__data_anchors_out),
.outs_ready (constant22_outs_ready__anchors_in),
.outs_valid (constant22_outs_valid__anchors_out),
.rst (rst)
);

extsi #(.INPUT_TYPE(2), .OUTPUT_TYPE(7)) extsi38(
.clk (clk),
.ins (constant22_outs__data_anchors_in),
.ins_ready (constant22_outs_ready__anchors_out),
.ins_valid (constant22_outs_valid__anchors_in),
.outs (extsi38_outs__data_anchors_out),
.outs_ready (extsi38_outs_ready__anchors_in),
.outs_valid (extsi38_outs_valid__anchors_out),
.rst (rst)
);

mc_store #(.DATA_TYPE(32), .ADDR_TYPE(32)) mc_store0(
.addrIn (extsi36_outs__data_anchors_in),
.addrIn_ready (extsi36_outs_ready__anchors_out),
.addrIn_valid (extsi36_outs_valid__anchors_in),
.addrOut (mc_store0_addrOut),
.addrOut_ready (mc_store0_addrOut_ready),
.addrOut_valid (mc_store0_addrOut_valid),
.clk (clk),
.dataIn (fork15_outs_1__data_anchors_in),
.dataIn_ready (fork15_outs_1_ready__anchors_out),
.dataIn_valid (fork15_outs_1_valid__anchors_in),
.dataToMem (mc_store0_dataToMem),
.dataToMem_ready (mc_store0_dataToMem_ready),
.dataToMem_valid (mc_store0_dataToMem_valid),
.rst (rst)
);

addi #(.DATA_TYPE(7)) addi14(
.clk (clk),
.lhs (extsi35_outs__data_anchors_in),
.lhs_ready (extsi35_outs_ready__anchors_out),
.lhs_valid (extsi35_outs_valid__anchors_in),
.result (addi14_result__data_anchors_out),
.result_ready (addi14_result_ready__anchors_in),
.result_valid (addi14_result_valid__anchors_out),
.rhs (extsi38_outs__data_anchors_in),
.rhs_ready (extsi38_outs_ready__anchors_out),
.rhs_valid (extsi38_outs_valid__anchors_in),
.rst (rst)
);

fork_type #(.SIZE(2), .DATA_TYPE(7)) fork17(
.clk (clk),
.ins (addi14_result__data_anchors_in),
.ins_ready (addi14_result_ready__anchors_out),
.ins_valid (addi14_result_valid__anchors_in),
.outs ({fork17_outs_1__data_anchors_out, fork17_outs_0__data_anchors_out}),
.outs_ready ({fork17_outs_1_ready__anchors_in, fork17_outs_0_ready__anchors_in}),
.outs_valid ({fork17_outs_1_valid__anchors_out, fork17_outs_0_valid__anchors_out}),
.rst (rst)
);

trunci #(.INPUT_TYPE(7), .OUTPUT_TYPE(6)) trunci2(
.clk (clk),
.ins (fork17_outs_0__data_anchors_in),
.ins_ready (fork17_outs_0_ready__anchors_out),
.ins_valid (fork17_outs_0_valid__anchors_in),
.outs (trunci2_outs__data_anchors_out),
.outs_ready (trunci2_outs_ready__anchors_in),
.outs_valid (trunci2_outs_valid__anchors_out),
.rst (rst)
);

handshake_cmpi_1 #(.DATA_TYPE(7)) cmpi5(
.clk (clk),
.lhs (fork17_outs_1__data_anchors_in),
.lhs_ready (fork17_outs_1_ready__anchors_out),
.lhs_valid (fork17_outs_1_valid__anchors_in),
.result (cmpi5_result__data_anchors_out),
.result_ready (cmpi5_result_ready__anchors_in),
.result_valid (cmpi5_result_valid__anchors_out),
.rhs (extsi37_outs__data_anchors_in),
.rhs_ready (extsi37_outs_ready__anchors_out),
.rhs_valid (extsi37_outs_valid__anchors_in),
.rst (rst)
);

fork_type #(.SIZE(3), .DATA_TYPE(1)) fork18(
.clk (clk),
.ins (cmpi5_result__data_anchors_in),
.ins_ready (cmpi5_result_ready__anchors_out),
.ins_valid (cmpi5_result_valid__anchors_in),
.outs ({fork18_outs_2__data_anchors_out, fork18_outs_1__data_anchors_out, fork18_outs_0__data_anchors_out}),
.outs_ready ({fork18_outs_2_ready__anchors_in, fork18_outs_1_ready__anchors_in, fork18_outs_0_ready__anchors_in}),
.outs_valid ({fork18_outs_2_valid__anchors_out, fork18_outs_1_valid__anchors_out, fork18_outs_0_valid__anchors_out}),
.rst (rst)
);

cond_br #(.DATA_TYPE(6)) cond_br17(
.clk (clk),
.condition (fork18_outs_0__data_anchors_in),
.condition_ready (fork18_outs_0_ready__anchors_out),
.condition_valid (fork18_outs_0_valid__anchors_in),
.data (trunci2_outs__data_anchors_in),
.data_ready (trunci2_outs_ready__anchors_out),
.data_valid (trunci2_outs_valid__anchors_in),
.falseOut (cond_br17_falseOut__data_anchors_out),
.falseOut_ready (cond_br17_falseOut_ready__anchors_in),
.falseOut_valid (cond_br17_falseOut_valid__anchors_out),
.rst (rst),
.trueOut (cond_br17_trueOut__data_anchors_out),
.trueOut_ready (cond_br17_trueOut_ready__anchors_in),
.trueOut_valid (cond_br17_trueOut_valid__anchors_out)
);

sink #(.DATA_TYPE(6)) sink4(
.clk (clk),
.ins (cond_br17_falseOut__data_anchors_in),
.ins_ready (cond_br17_falseOut_ready__anchors_out),
.ins_valid (cond_br17_falseOut_valid__anchors_in),
.rst (rst)
);

cond_br_dataless cond_br13(
.clk (clk),
.condition (fork18_outs_1__data_anchors_in),
.condition_ready (fork18_outs_1_ready__anchors_out),
.condition_valid (fork18_outs_1_valid__anchors_in),
.data_ready (fork16_outs_1_ready__anchors_out),
.data_valid (fork16_outs_1_valid__anchors_in),
.falseOut_ready (cond_br13_falseOut_ready__anchors_in),
.falseOut_valid (cond_br13_falseOut_valid__anchors_out),
.rst (rst),
.trueOut_ready (cond_br13_trueOut_ready__anchors_in),
.trueOut_valid (cond_br13_trueOut_valid__anchors_out)
);

cond_br #(.DATA_TYPE(32)) cond_br14(
.clk (clk),
.condition (fork18_outs_2__data_anchors_in),
.condition_ready (fork18_outs_2_ready__anchors_out),
.condition_valid (fork18_outs_2_valid__anchors_in),
.data (fork15_outs_0__data_anchors_in),
.data_ready (fork15_outs_0_ready__anchors_out),
.data_valid (fork15_outs_0_valid__anchors_in),
.falseOut (cond_br14_falseOut__data_anchors_out),
.falseOut_ready (cond_br14_falseOut_ready__anchors_in),
.falseOut_valid (cond_br14_falseOut_valid__anchors_out),
.rst (rst),
.trueOut (cond_br14_trueOut__data_anchors_out),
.trueOut_ready (cond_br14_trueOut_ready__anchors_in),
.trueOut_valid (cond_br14_trueOut_valid__anchors_out)
);

sink #(.DATA_TYPE(32)) sink5(
.clk (clk),
.ins (cond_br14_trueOut__data_anchors_in),
.ins_ready (cond_br14_trueOut_ready__anchors_out),
.ins_valid (cond_br14_trueOut_valid__anchors_in),
.rst (rst)
);

fork_dataless #(.SIZE(3)) fork19(
.clk (clk),
.ins_ready (cond_br13_falseOut_ready__anchors_out),
.ins_valid (cond_br13_falseOut_valid__anchors_in),
.outs_ready ({fork19_outs_2_ready__anchors_in, fork19_outs_1_ready__anchors_in, fork19_outs_0_ready__anchors_in}),
.outs_valid ({fork19_outs_2_valid__anchors_out, fork19_outs_1_valid__anchors_out, fork19_outs_0_valid__anchors_out}),
.rst (rst)
);

endmodule
